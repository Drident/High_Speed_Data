library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package nxPackage is

-- FAMILY

constant NX_SYMBOL : string := "NG_M";
constant NX_FAMILY : string := "NG_MEDIUM";

-- IOM

constant IOM_LINK_DES_CHAIN_IN          : integer := 0;
constant IOM_LINK_SER_FCK_FABRIC        : integer := 1;
constant IOM_LINK_CTCK_FABRIC           : integer := 2;
constant IOM_LINK_SPW_TX_SO             : integer := 3;
constant IOM_LINK_DES_FCK_FABRIC        : integer := 4;
constant IOM_LINK_SPW_TX_OUT_CONFIG     : integer := 5;
constant IOM_LINK_SER_WPTR              : integer := 6;
constant IOM_LINK_SER_SCK_IOM           : integer := 7;
constant IOM_LINK_FZ                    : integer := 8;
constant IOM_LINK_SPW_RX_RCK            : integer := 9;
constant IOM_LINK_SER_CHAIN_IN          : integer := 10;
constant IOM_LINK_SER_RPTR              : integer := 11;
constant IOM_LINK_DES_SCK_IOM           : integer := 12;
constant IOM_LINK_DELAY_VALUE_IN_LAST   : integer := 13;
constant IOM_LINK_DELAY_VALUE_IN_FIRST  : integer := 18;
constant IOM_LINK_SPW_RX_DI             : integer := 19;
constant IOM_LINK_DCK                   : integer := 20;
constant IOM_LINK_DWR                   : integer := 21;
constant IOM_LINK_DES_RPTR              : integer := 22;
constant IOM_LINK_SER_SCK_FABRIC        : integer := 23;
constant IOM_LINK_DELAY_SELECT_LAST     : integer := 24;
constant IOM_LINK_DELAY_SELECT_FIRST    : integer := 25;
constant IOM_LINK_SPW_RX_IN_CONFIG      : integer := 26;
constant IOM_LINK_DES_WPTR              : integer := 27;
constant IOM_LINK_DES_SCK_FABRIC        : integer := 28;
constant IOM_LINK_SPW_TX_DO             : integer := 29;
constant IOM_LINK_SPW_RX_DATA           : integer := 30;
constant IOM_LINK_DES_CHAIN_OUT         : integer := 31;
constant IOM_LINK_DELAY_VALUE_OUT_LAST  : integer := 32;
constant IOM_LINK_DELAY_VALUE_OUT_FIRST : integer := 37;
constant IOM_LINK_FLD                   : integer := 38;
constant IOM_LINK_SER_CHAIN_OUT         : integer := 39;
constant IOM_LINK_FLG                   : integer := 40;
constant IOM_LINK_PAD_SYSCLK            : integer := 41;
constant IOM_LINK_SIZE                  : integer := 42;
constant IOM_LINK_OUTPUT_MAX            : integer := 28;

-- HSSL

constant CRX_LINK_SIZE                  : integer := 10;

constant CTX_LINK_SIZE                  : integer := 20;

component NX_CDC_L is
generic (
    mode : bit := '0';
    rck_edge : bit := '0';
    wck_edge : bit := '0'
);
port (
    CK	: in std_logic := '0';
    RI1	: in std_logic := '0';
    RI2	: in std_logic := '0';
    RI3	: in std_logic := '0';
    RI4	: in std_logic := '0';
    RI5	: in std_logic := '0';
    RI6	: in std_logic := '0';
    RO1	: out std_logic := '0';
    RO2	: out std_logic := '0';
    RO3	: out std_logic := '0';
    RO4	: out std_logic := '0';
    RO5	: out std_logic := '0';
    RO6	: out std_logic := '0';
    WI1	: in std_logic := '0';
    WI2	: in std_logic := '0';
    WI3	: in std_logic := '0';
    WI4	: in std_logic := '0';
    WI5	: in std_logic := '0';
    WI6	: in std_logic := '0';
    WO1	: out std_logic := '0';
    WO2	: out std_logic := '0';
    WO3	: out std_logic := '0';
    WO4	: out std_logic := '0';
    WO5	: out std_logic := '0';
    WO6	: out std_logic := '0'
);
end component NX_CDC_L;

component NX_FIFO_CDC_L is
generic (
    mode : bit := '1'
);
port (
    XRCK	: in std_logic := '0';
    XWCK	: in std_logic := '0';
    XRI1	: in std_logic := '0';
    XRI2	: in std_logic := '0';
    XRI3	: in std_logic := '0';
    XRI4	: in std_logic := '0';
    XRI5	: in std_logic := '0';
    XRI6	: in std_logic := '0';
    XWI1	: in std_logic := '0';
    XWI2	: in std_logic := '0';
    XWI3	: in std_logic := '0';
    XWI4	: in std_logic := '0';
    XWI5	: in std_logic := '0';
    XWI6	: in std_logic := '0';
    RO1	: out std_logic := '0';
    RO2	: out std_logic := '0';
    RO3	: out std_logic := '0';
    RO4	: out std_logic := '0';
    RO5	: out std_logic := '0';
    RO6	: out std_logic := '0';
    WO1	: out std_logic := '0';
    WO2	: out std_logic := '0';
    WO3	: out std_logic := '0';
    WO4	: out std_logic := '0';
    WO5	: out std_logic := '0';
    WO6	: out std_logic := '0'
);
end component NX_FIFO_CDC_L;

component NX_DSPDPRAM_FULL_L is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    dsp0_clk_i	: in std_logic := '0';
    dsp0_rst_i	: in std_logic := '0';
    dsp0_rstz_i	: in std_logic := '0';
    dsp0_we_i	: in std_logic := '0';
    dsp0_cy_i	: in std_logic := '0';
    dsp0_a_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dsp0_b_i	: in std_logic_vector(17 downto 0) := (others => '0');
    dsp0_c_i	: in std_logic_vector(35 downto 0) := (others => '0');
    dsp0_d_i	: in std_logic_vector(17 downto 0) := (others => '0');

    dsp0_z_o	: out std_logic_vector(55 downto 0) := (others => '0');
    dsp0_cy_o	: out std_logic := '0';
    dsp0_cy36_o	: out std_logic := '0';
    dsp0_cy56_o	: out std_logic := '0';
    dsp0_ovf_o	: out std_logic := '0';

    dsp1_clk_i	: in std_logic := '0';
    dsp1_rst_i	: in std_logic := '0';
    dsp1_rstz_i	: in std_logic := '0';
    dsp1_we_i	: in std_logic := '0';
    dsp1_cy_i	: in std_logic := '0';
    dsp1_a_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dsp1_b_i	: in std_logic_vector(17 downto 0) := (others => '0');
    dsp1_c_i	: in std_logic_vector(35 downto 0) := (others => '0');
    dsp1_d_i	: in std_logic_vector(17 downto 0) := (others => '0');

    dsp1_z_o	: out std_logic_vector(55 downto 0) := (others => '0');
    dsp1_cy_o	: out std_logic := '0';
    dsp1_cy36_o	: out std_logic := '0';
    dsp1_cy56_o	: out std_logic := '0';
    dsp1_ovf_o	: out std_logic := '0';

    dsp_ca_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dsp_cb_i	: in std_logic_vector(17 downto 0) := (others => '0');
    dsp_cz_i	: in std_logic_vector(55 downto 0) := (others => '0');
    dsp_ccy_i	: in std_logic := '0';
    dsp_ca_o	: out std_logic_vector(23 downto 0) := (others => '0');
    dsp_cb_o	: out std_logic_vector(17 downto 0) := (others => '0');
    dsp_cz_o	: out std_logic_vector(55 downto 0) := (others => '0');
    dsp_ccy_o	: out std_logic := '0';


    dpram_clkmem0_i	: in std_logic := '0';
    dpram_clkmemclone0_i	: in std_logic := '0';
    dpram_clkmem90_0_i	: in std_logic := '0';
    dpram_clkreg0_i	: in std_logic := '0';
    dpram_rst0_i	: in std_logic := '0';
    dpram_cs0_i	: in std_logic := '0';
    dpram_we0_i	: in std_logic := '0';
    dpram_addr0_i	: in std_logic_vector(15 downto 0) := (others => '0');
    dpram_din0_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dpram_dout0_o	: out std_logic_vector(23 downto 0) := (others => '0');
    dpram_ecc_corrected0_o	: out std_logic := '0';
    dpram_ecc_uncorrected0_o	: out std_logic := '0';

    dpram_clkmem1_i	: in std_logic := '0';
    dpram_clkmemclone1_i	: in std_logic := '0';
    dpram_clkmem90_1_i	: in std_logic := '0';
    dpram_clkreg1_i	: in std_logic := '0';
    dpram_rst1_i	: in std_logic := '0';
    dpram_cs1_i	: in std_logic := '0';
    dpram_we1_i	: in std_logic := '0';
    dpram_addr1_i	: in std_logic_vector(15 downto 0) := (others => '0');
    dpram_din1_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dpram_dout1_o	: out std_logic_vector(23 downto 0) := (others => '0');
    dpram_ecc_corrected1_o	: out std_logic := '0';
    dpram_ecc_uncorrected1_o	: out std_logic := '0'
);
end component NX_DSPDPRAM_FULL_L;

component NX_DSP_L_BOX is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    A5	: in std_logic := '0';
    A6	: in std_logic := '0';
    A7	: in std_logic := '0';
    A8	: in std_logic := '0';
    A9	: in std_logic := '0';
    A10	: in std_logic := '0';
    A11	: in std_logic := '0';
    A12	: in std_logic := '0';
    A13	: in std_logic := '0';
    A14	: in std_logic := '0';
    A15	: in std_logic := '0';
    A16	: in std_logic := '0';
    A17	: in std_logic := '0';
    A18	: in std_logic := '0';
    A19	: in std_logic := '0';
    A20	: in std_logic := '0';
    A21	: in std_logic := '0';
    A22	: in std_logic := '0';
    A23	: in std_logic := '0';
    A24	: in std_logic := '0';

    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    B5	: in std_logic := '0';
    B6	: in std_logic := '0';
    B7	: in std_logic := '0';
    B8	: in std_logic := '0';
    B9	: in std_logic := '0';
    B10	: in std_logic := '0';
    B11	: in std_logic := '0';
    B12	: in std_logic := '0';
    B13	: in std_logic := '0';
    B14	: in std_logic := '0';
    B15	: in std_logic := '0';
    B16	: in std_logic := '0';
    B17	: in std_logic := '0';
    B18	: in std_logic := '0';

    C1	: in std_logic := '0';
    C2	: in std_logic := '0';
    C3	: in std_logic := '0';
    C4	: in std_logic := '0';
    C5	: in std_logic := '0';
    C6	: in std_logic := '0';
    C7	: in std_logic := '0';
    C8	: in std_logic := '0';
    C9	: in std_logic := '0';
    C10	: in std_logic := '0';
    C11	: in std_logic := '0';
    C12	: in std_logic := '0';
    C13	: in std_logic := '0';
    C14	: in std_logic := '0';
    C15	: in std_logic := '0';
    C16	: in std_logic := '0';
    C17	: in std_logic := '0';
    C18	: in std_logic := '0';
    C19	: in std_logic := '0';
    C20	: in std_logic := '0';
    C21	: in std_logic := '0';
    C22	: in std_logic := '0';
    C23	: in std_logic := '0';
    C24	: in std_logic := '0';
    C25	: in std_logic := '0';
    C26	: in std_logic := '0';
    C27	: in std_logic := '0';
    C28	: in std_logic := '0';
    C29	: in std_logic := '0';
    C30	: in std_logic := '0';
    C31	: in std_logic := '0';
    C32	: in std_logic := '0';
    C33	: in std_logic := '0';
    C34	: in std_logic := '0';
    C35	: in std_logic := '0';
    C36	: in std_logic := '0';

    CAI1	: in std_logic := '0';
    CAI2	: in std_logic := '0';
    CAI3	: in std_logic := '0';
    CAI4	: in std_logic := '0';
    CAI5	: in std_logic := '0';
    CAI6	: in std_logic := '0';
    CAI7	: in std_logic := '0';
    CAI8	: in std_logic := '0';
    CAI9	: in std_logic := '0';
    CAI10	: in std_logic := '0';
    CAI11	: in std_logic := '0';
    CAI12	: in std_logic := '0';
    CAI13	: in std_logic := '0';
    CAI14	: in std_logic := '0';
    CAI15	: in std_logic := '0';
    CAI16	: in std_logic := '0';
    CAI17	: in std_logic := '0';
    CAI18	: in std_logic := '0';
    CAI19	: in std_logic := '0';
    CAI20	: in std_logic := '0';
    CAI21	: in std_logic := '0';
    CAI22	: in std_logic := '0';
    CAI23	: in std_logic := '0';
    CAI24	: in std_logic := '0';

    CAO1	: out std_logic := '0';
    CAO2	: out std_logic := '0';
    CAO3	: out std_logic := '0';
    CAO4	: out std_logic := '0';
    CAO5	: out std_logic := '0';
    CAO6	: out std_logic := '0';
    CAO7	: out std_logic := '0';
    CAO8	: out std_logic := '0';
    CAO9	: out std_logic := '0';
    CAO10	: out std_logic := '0';
    CAO11	: out std_logic := '0';
    CAO12	: out std_logic := '0';
    CAO13	: out std_logic := '0';
    CAO14	: out std_logic := '0';
    CAO15	: out std_logic := '0';
    CAO16	: out std_logic := '0';
    CAO17	: out std_logic := '0';
    CAO18	: out std_logic := '0';
    CAO19	: out std_logic := '0';
    CAO20	: out std_logic := '0';
    CAO21	: out std_logic := '0';
    CAO22	: out std_logic := '0';
    CAO23	: out std_logic := '0';
    CAO24	: out std_logic := '0';

    CBI1	: in std_logic := '0';
    CBI2	: in std_logic := '0';
    CBI3	: in std_logic := '0';
    CBI4	: in std_logic := '0';
    CBI5	: in std_logic := '0';
    CBI6	: in std_logic := '0';
    CBI7	: in std_logic := '0';
    CBI8	: in std_logic := '0';
    CBI9	: in std_logic := '0';
    CBI10	: in std_logic := '0';
    CBI11	: in std_logic := '0';
    CBI12	: in std_logic := '0';
    CBI13	: in std_logic := '0';
    CBI14	: in std_logic := '0';
    CBI15	: in std_logic := '0';
    CBI16	: in std_logic := '0';
    CBI17	: in std_logic := '0';
    CBI18	: in std_logic := '0';

    CBO1	: out std_logic := '0';
    CBO2	: out std_logic := '0';
    CBO3	: out std_logic := '0';
    CBO4	: out std_logic := '0';
    CBO5	: out std_logic := '0';
    CBO6	: out std_logic := '0';
    CBO7	: out std_logic := '0';
    CBO8	: out std_logic := '0';
    CBO9	: out std_logic := '0';
    CBO10	: out std_logic := '0';
    CBO11	: out std_logic := '0';
    CBO12	: out std_logic := '0';
    CBO13	: out std_logic := '0';
    CBO14	: out std_logic := '0';
    CBO15	: out std_logic := '0';
    CBO16	: out std_logic := '0';
    CBO17	: out std_logic := '0';
    CBO18	: out std_logic := '0';

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO	: out std_logic := '0';
    CO37	: out std_logic := '0';
    CO57	: out std_logic := '0';

    CZI1	: in std_logic := '0';
    CZI2	: in std_logic := '0';
    CZI3	: in std_logic := '0';
    CZI4	: in std_logic := '0';
    CZI5	: in std_logic := '0';
    CZI6	: in std_logic := '0';
    CZI7	: in std_logic := '0';
    CZI8	: in std_logic := '0';
    CZI9	: in std_logic := '0';
    CZI10	: in std_logic := '0';
    CZI11	: in std_logic := '0';
    CZI12	: in std_logic := '0';
    CZI13	: in std_logic := '0';
    CZI14	: in std_logic := '0';
    CZI15	: in std_logic := '0';
    CZI16	: in std_logic := '0';
    CZI17	: in std_logic := '0';
    CZI18	: in std_logic := '0';
    CZI19	: in std_logic := '0';
    CZI20	: in std_logic := '0';
    CZI21	: in std_logic := '0';
    CZI22	: in std_logic := '0';
    CZI23	: in std_logic := '0';
    CZI24	: in std_logic := '0';
    CZI25	: in std_logic := '0';
    CZI26	: in std_logic := '0';
    CZI27	: in std_logic := '0';
    CZI28	: in std_logic := '0';
    CZI29	: in std_logic := '0';
    CZI30	: in std_logic := '0';
    CZI31	: in std_logic := '0';
    CZI32	: in std_logic := '0';
    CZI33	: in std_logic := '0';
    CZI34	: in std_logic := '0';
    CZI35	: in std_logic := '0';
    CZI36	: in std_logic := '0';
    CZI37	: in std_logic := '0';
    CZI38	: in std_logic := '0';
    CZI39	: in std_logic := '0';
    CZI40	: in std_logic := '0';
    CZI41	: in std_logic := '0';
    CZI42	: in std_logic := '0';
    CZI43	: in std_logic := '0';
    CZI44	: in std_logic := '0';
    CZI45	: in std_logic := '0';
    CZI46	: in std_logic := '0';
    CZI47	: in std_logic := '0';
    CZI48	: in std_logic := '0';
    CZI49	: in std_logic := '0';
    CZI50	: in std_logic := '0';
    CZI51	: in std_logic := '0';
    CZI52	: in std_logic := '0';
    CZI53	: in std_logic := '0';
    CZI54	: in std_logic := '0';
    CZI55	: in std_logic := '0';
    CZI56	: in std_logic := '0';

    CZO1	: out std_logic := '0';
    CZO2	: out std_logic := '0';
    CZO3	: out std_logic := '0';
    CZO4	: out std_logic := '0';
    CZO5	: out std_logic := '0';
    CZO6	: out std_logic := '0';
    CZO7	: out std_logic := '0';
    CZO8	: out std_logic := '0';
    CZO9	: out std_logic := '0';
    CZO10	: out std_logic := '0';
    CZO11	: out std_logic := '0';
    CZO12	: out std_logic := '0';
    CZO13	: out std_logic := '0';
    CZO14	: out std_logic := '0';
    CZO15	: out std_logic := '0';
    CZO16	: out std_logic := '0';
    CZO17	: out std_logic := '0';
    CZO18	: out std_logic := '0';
    CZO19	: out std_logic := '0';
    CZO20	: out std_logic := '0';
    CZO21	: out std_logic := '0';
    CZO22	: out std_logic := '0';
    CZO23	: out std_logic := '0';
    CZO24	: out std_logic := '0';
    CZO25	: out std_logic := '0';
    CZO26	: out std_logic := '0';
    CZO27	: out std_logic := '0';
    CZO28	: out std_logic := '0';
    CZO29	: out std_logic := '0';
    CZO30	: out std_logic := '0';
    CZO31	: out std_logic := '0';
    CZO32	: out std_logic := '0';
    CZO33	: out std_logic := '0';
    CZO34	: out std_logic := '0';
    CZO35	: out std_logic := '0';
    CZO36	: out std_logic := '0';
    CZO37	: out std_logic := '0';
    CZO38	: out std_logic := '0';
    CZO39	: out std_logic := '0';
    CZO40	: out std_logic := '0';
    CZO41	: out std_logic := '0';
    CZO42	: out std_logic := '0';
    CZO43	: out std_logic := '0';
    CZO44	: out std_logic := '0';
    CZO45	: out std_logic := '0';
    CZO46	: out std_logic := '0';
    CZO47	: out std_logic := '0';
    CZO48	: out std_logic := '0';
    CZO49	: out std_logic := '0';
    CZO50	: out std_logic := '0';
    CZO51	: out std_logic := '0';
    CZO52	: out std_logic := '0';
    CZO53	: out std_logic := '0';
    CZO54	: out std_logic := '0';
    CZO55	: out std_logic := '0';
    CZO56	: out std_logic := '0';

    D1	: in std_logic := '0';
    D2	: in std_logic := '0';
    D3	: in std_logic := '0';
    D4	: in std_logic := '0';
    D5	: in std_logic := '0';
    D6	: in std_logic := '0';
    D7	: in std_logic := '0';
    D8	: in std_logic := '0';
    D9	: in std_logic := '0';
    D10	: in std_logic := '0';
    D11	: in std_logic := '0';
    D12	: in std_logic := '0';
    D13	: in std_logic := '0';
    D14	: in std_logic := '0';
    D15	: in std_logic := '0';
    D16	: in std_logic := '0';
    D17	: in std_logic := '0';
    D18	: in std_logic := '0';

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';

    Z1	: out std_logic := '0';
    Z2	: out std_logic := '0';
    Z3	: out std_logic := '0';
    Z4	: out std_logic := '0';
    Z5	: out std_logic := '0';
    Z6	: out std_logic := '0';
    Z7	: out std_logic := '0';
    Z8	: out std_logic := '0';
    Z9	: out std_logic := '0';
    Z10	: out std_logic := '0';
    Z11	: out std_logic := '0';
    Z12	: out std_logic := '0';
    Z13	: out std_logic := '0';
    Z14	: out std_logic := '0';
    Z15	: out std_logic := '0';
    Z16	: out std_logic := '0';
    Z17	: out std_logic := '0';
    Z18	: out std_logic := '0';
    Z19	: out std_logic := '0';
    Z20	: out std_logic := '0';
    Z21	: out std_logic := '0';
    Z22	: out std_logic := '0';
    Z23	: out std_logic := '0';
    Z24	: out std_logic := '0';
    Z25	: out std_logic := '0';
    Z26	: out std_logic := '0';
    Z27	: out std_logic := '0';
    Z28	: out std_logic := '0';
    Z29	: out std_logic := '0';
    Z30	: out std_logic := '0';
    Z31	: out std_logic := '0';
    Z32	: out std_logic := '0';
    Z33	: out std_logic := '0';
    Z34	: out std_logic := '0';
    Z35	: out std_logic := '0';
    Z36	: out std_logic := '0';
    Z37	: out std_logic := '0';
    Z38	: out std_logic := '0';
    Z39	: out std_logic := '0';
    Z40	: out std_logic := '0';
    Z41	: out std_logic := '0';
    Z42	: out std_logic := '0';
    Z43	: out std_logic := '0';
    Z44	: out std_logic := '0';
    Z45	: out std_logic := '0';
    Z46	: out std_logic := '0';
    Z47	: out std_logic := '0';
    Z48	: out std_logic := '0';
    Z49	: out std_logic := '0';
    Z50	: out std_logic := '0';
    Z51	: out std_logic := '0';
    Z52	: out std_logic := '0';
    Z53	: out std_logic := '0';
    Z54	: out std_logic := '0';
    Z55	: out std_logic := '0';
    Z56	: out std_logic := '0'
);
end component NX_DSP_L_BOX;

component NX_RAM_L_BOX is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    ACK	: in std_logic := '0';
    ACKC	: in std_logic := '0';
    ACKD	: in std_logic := '0';
    ACKR	: in std_logic := '0';
    BCK	: in std_logic := '0';
    BCKC	: in std_logic := '0';
    BCKD	: in std_logic := '0';
    BCKR	: in std_logic := '0';

    AI1	: in std_logic := '0';
    AI2	: in std_logic := '0';
    AI3	: in std_logic := '0';
    AI4	: in std_logic := '0';
    AI5	: in std_logic := '0';
    AI6	: in std_logic := '0';
    AI7	: in std_logic := '0';
    AI8	: in std_logic := '0';
    AI9	: in std_logic := '0';
    AI10	: in std_logic := '0';
    AI11	: in std_logic := '0';
    AI12	: in std_logic := '0';
    AI13	: in std_logic := '0';
    AI14	: in std_logic := '0';
    AI15	: in std_logic := '0';
    AI16	: in std_logic := '0';

    AI17	: in std_logic := '0';
    AI18	: in std_logic := '0';
    AI19	: in std_logic := '0';
    AI20	: in std_logic := '0';
    AI21	: in std_logic := '0';
    AI22	: in std_logic := '0';
    AI23	: in std_logic := '0';
    AI24	: in std_logic := '0';

    BI1	: in std_logic := '0';
    BI2	: in std_logic := '0';
    BI3	: in std_logic := '0';
    BI4	: in std_logic := '0';
    BI5	: in std_logic := '0';
    BI6	: in std_logic := '0';
    BI7	: in std_logic := '0';
    BI8	: in std_logic := '0';
    BI9	: in std_logic := '0';
    BI10	: in std_logic := '0';
    BI11	: in std_logic := '0';
    BI12	: in std_logic := '0';
    BI13	: in std_logic := '0';
    BI14	: in std_logic := '0';
    BI15	: in std_logic := '0';
    BI16	: in std_logic := '0';

    BI17	: in std_logic := '0';
    BI18	: in std_logic := '0';
    BI19	: in std_logic := '0';
    BI20	: in std_logic := '0';
    BI21	: in std_logic := '0';
    BI22	: in std_logic := '0';
    BI23	: in std_logic := '0';
    BI24	: in std_logic := '0';

    ACOR	: out std_logic := '0';
    AERR	: out std_logic := '0';
    BCOR	: out std_logic := '0';
    BERR	: out std_logic := '0';

    AO1	: out std_logic := '0';
    AO2	: out std_logic := '0';
    AO3	: out std_logic := '0';
    AO4	: out std_logic := '0';
    AO5	: out std_logic := '0';
    AO6	: out std_logic := '0';
    AO7	: out std_logic := '0';
    AO8	: out std_logic := '0';
    AO9	: out std_logic := '0';
    AO10	: out std_logic := '0';
    AO11	: out std_logic := '0';
    AO12	: out std_logic := '0';
    AO13	: out std_logic := '0';
    AO14	: out std_logic := '0';
    AO15	: out std_logic := '0';
    AO16	: out std_logic := '0';

    AO17	: out std_logic := '0';
    AO18	: out std_logic := '0';
    AO19	: out std_logic := '0';
    AO20	: out std_logic := '0';
    AO21	: out std_logic := '0';
    AO22	: out std_logic := '0';
    AO23	: out std_logic := '0';
    AO24	: out std_logic := '0';

    BO1	: out std_logic := '0';
    BO2	: out std_logic := '0';
    BO3	: out std_logic := '0';
    BO4	: out std_logic := '0';
    BO5	: out std_logic := '0';
    BO6	: out std_logic := '0';
    BO7	: out std_logic := '0';
    BO8	: out std_logic := '0';
    BO9	: out std_logic := '0';
    BO10	: out std_logic := '0';
    BO11	: out std_logic := '0';
    BO12	: out std_logic := '0';
    BO13	: out std_logic := '0';
    BO14	: out std_logic := '0';
    BO15	: out std_logic := '0';
    BO16	: out std_logic := '0';

    BO17	: out std_logic := '0';
    BO18	: out std_logic := '0';
    BO19	: out std_logic := '0';
    BO20	: out std_logic := '0';
    BO21	: out std_logic := '0';
    BO22	: out std_logic := '0';
    BO23	: out std_logic := '0';
    BO24	: out std_logic := '0';

    AA1	: in std_logic := '0';
    AA2	: in std_logic := '0';
    AA3	: in std_logic := '0';
    AA4	: in std_logic := '0';
    AA5	: in std_logic := '0';
    AA6	: in std_logic := '0';

    AA7	: in std_logic := '0';
    AA8	: in std_logic := '0';
    AA9	: in std_logic := '0';
    AA10	: in std_logic := '0';
    AA11	: in std_logic := '0';
    AA12	: in std_logic := '0';
    AA13	: in std_logic := '0';
    AA14	: in std_logic := '0';
    AA15	: in std_logic := '0';
    AA16	: in std_logic := '0';

    ACS	: in std_logic := '0';
    AWE	: in std_logic := '0';
    AR	: in std_logic := '0';

    BA1	: in std_logic := '0';
    BA2	: in std_logic := '0';
    BA3	: in std_logic := '0';
    BA4	: in std_logic := '0';
    BA5	: in std_logic := '0';
    BA6	: in std_logic := '0';

    BA7	: in std_logic := '0';
    BA8	: in std_logic := '0';
    BA9	: in std_logic := '0';
    BA10	: in std_logic := '0';
    BA11	: in std_logic := '0';
    BA12	: in std_logic := '0';
    BA13	: in std_logic := '0';
    BA14	: in std_logic := '0';
    BA15	: in std_logic := '0';
    BA16	: in std_logic := '0';

    BCS	: in std_logic := '0';
    BWE	: in std_logic := '0';
    BR	: in std_logic := '0'
);
end component NX_RAM_L_BOX;

component NX_DSP_L is
generic (
    std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";   -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";    -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";          -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                 -- ALU
);
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    A5	: in std_logic := '0';
    A6	: in std_logic := '0';
    A7	: in std_logic := '0';
    A8	: in std_logic := '0';
    A9	: in std_logic := '0';
    A10	: in std_logic := '0';
    A11	: in std_logic := '0';
    A12	: in std_logic := '0';
    A13	: in std_logic := '0';
    A14	: in std_logic := '0';
    A15	: in std_logic := '0';
    A16	: in std_logic := '0';
    A17	: in std_logic := '0';
    A18	: in std_logic := '0';
    A19	: in std_logic := '0';
    A20	: in std_logic := '0';
    A21	: in std_logic := '0';
    A22	: in std_logic := '0';
    A23	: in std_logic := '0';
    A24	: in std_logic := '0';

    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    B5	: in std_logic := '0';
    B6	: in std_logic := '0';
    B7	: in std_logic := '0';
    B8	: in std_logic := '0';
    B9	: in std_logic := '0';
    B10	: in std_logic := '0';
    B11	: in std_logic := '0';
    B12	: in std_logic := '0';
    B13	: in std_logic := '0';
    B14	: in std_logic := '0';
    B15	: in std_logic := '0';
    B16	: in std_logic := '0';
    B17	: in std_logic := '0';
    B18	: in std_logic := '0';

    C1	: in std_logic := '0';
    C2	: in std_logic := '0';
    C3	: in std_logic := '0';
    C4	: in std_logic := '0';
    C5	: in std_logic := '0';
    C6	: in std_logic := '0';
    C7	: in std_logic := '0';
    C8	: in std_logic := '0';
    C9	: in std_logic := '0';
    C10	: in std_logic := '0';
    C11	: in std_logic := '0';
    C12	: in std_logic := '0';
    C13	: in std_logic := '0';
    C14	: in std_logic := '0';
    C15	: in std_logic := '0';
    C16	: in std_logic := '0';
    C17	: in std_logic := '0';
    C18	: in std_logic := '0';
    C19	: in std_logic := '0';
    C20	: in std_logic := '0';
    C21	: in std_logic := '0';
    C22	: in std_logic := '0';
    C23	: in std_logic := '0';
    C24	: in std_logic := '0';
    C25	: in std_logic := '0';
    C26	: in std_logic := '0';
    C27	: in std_logic := '0';
    C28	: in std_logic := '0';
    C29	: in std_logic := '0';
    C30	: in std_logic := '0';
    C31	: in std_logic := '0';
    C32	: in std_logic := '0';
    C33	: in std_logic := '0';
    C34	: in std_logic := '0';
    C35	: in std_logic := '0';
    C36	: in std_logic := '0';

    CAI1	: in std_logic := '0';
    CAI2	: in std_logic := '0';
    CAI3	: in std_logic := '0';
    CAI4	: in std_logic := '0';
    CAI5	: in std_logic := '0';
    CAI6	: in std_logic := '0';
    CAI7	: in std_logic := '0';
    CAI8	: in std_logic := '0';
    CAI9	: in std_logic := '0';
    CAI10	: in std_logic := '0';
    CAI11	: in std_logic := '0';
    CAI12	: in std_logic := '0';
    CAI13	: in std_logic := '0';
    CAI14	: in std_logic := '0';
    CAI15	: in std_logic := '0';
    CAI16	: in std_logic := '0';
    CAI17	: in std_logic := '0';
    CAI18	: in std_logic := '0';
    CAI19	: in std_logic := '0';
    CAI20	: in std_logic := '0';
    CAI21	: in std_logic := '0';
    CAI22	: in std_logic := '0';
    CAI23	: in std_logic := '0';
    CAI24	: in std_logic := '0';

    CAO1	: out std_logic := '0';
    CAO2	: out std_logic := '0';
    CAO3	: out std_logic := '0';
    CAO4	: out std_logic := '0';
    CAO5	: out std_logic := '0';
    CAO6	: out std_logic := '0';
    CAO7	: out std_logic := '0';
    CAO8	: out std_logic := '0';
    CAO9	: out std_logic := '0';
    CAO10	: out std_logic := '0';
    CAO11	: out std_logic := '0';
    CAO12	: out std_logic := '0';
    CAO13	: out std_logic := '0';
    CAO14	: out std_logic := '0';
    CAO15	: out std_logic := '0';
    CAO16	: out std_logic := '0';
    CAO17	: out std_logic := '0';
    CAO18	: out std_logic := '0';
    CAO19	: out std_logic := '0';
    CAO20	: out std_logic := '0';
    CAO21	: out std_logic := '0';
    CAO22	: out std_logic := '0';
    CAO23	: out std_logic := '0';
    CAO24	: out std_logic := '0';

    CBI1	: in std_logic := '0';
    CBI2	: in std_logic := '0';
    CBI3	: in std_logic := '0';
    CBI4	: in std_logic := '0';
    CBI5	: in std_logic := '0';
    CBI6	: in std_logic := '0';
    CBI7	: in std_logic := '0';
    CBI8	: in std_logic := '0';
    CBI9	: in std_logic := '0';
    CBI10	: in std_logic := '0';
    CBI11	: in std_logic := '0';
    CBI12	: in std_logic := '0';
    CBI13	: in std_logic := '0';
    CBI14	: in std_logic := '0';
    CBI15	: in std_logic := '0';
    CBI16	: in std_logic := '0';
    CBI17	: in std_logic := '0';
    CBI18	: in std_logic := '0';

    CBO1	: out std_logic := '0';
    CBO2	: out std_logic := '0';
    CBO3	: out std_logic := '0';
    CBO4	: out std_logic := '0';
    CBO5	: out std_logic := '0';
    CBO6	: out std_logic := '0';
    CBO7	: out std_logic := '0';
    CBO8	: out std_logic := '0';
    CBO9	: out std_logic := '0';
    CBO10	: out std_logic := '0';
    CBO11	: out std_logic := '0';
    CBO12	: out std_logic := '0';
    CBO13	: out std_logic := '0';
    CBO14	: out std_logic := '0';
    CBO15	: out std_logic := '0';
    CBO16	: out std_logic := '0';
    CBO17	: out std_logic := '0';
    CBO18	: out std_logic := '0';

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO	: out std_logic := '0';
    CO37	: out std_logic := '0';
    CO57	: out std_logic := '0';

    CZI1	: in std_logic := '0';
    CZI2	: in std_logic := '0';
    CZI3	: in std_logic := '0';
    CZI4	: in std_logic := '0';
    CZI5	: in std_logic := '0';
    CZI6	: in std_logic := '0';
    CZI7	: in std_logic := '0';
    CZI8	: in std_logic := '0';
    CZI9	: in std_logic := '0';
    CZI10	: in std_logic := '0';
    CZI11	: in std_logic := '0';
    CZI12	: in std_logic := '0';
    CZI13	: in std_logic := '0';
    CZI14	: in std_logic := '0';
    CZI15	: in std_logic := '0';
    CZI16	: in std_logic := '0';
    CZI17	: in std_logic := '0';
    CZI18	: in std_logic := '0';
    CZI19	: in std_logic := '0';
    CZI20	: in std_logic := '0';
    CZI21	: in std_logic := '0';
    CZI22	: in std_logic := '0';
    CZI23	: in std_logic := '0';
    CZI24	: in std_logic := '0';
    CZI25	: in std_logic := '0';
    CZI26	: in std_logic := '0';
    CZI27	: in std_logic := '0';
    CZI28	: in std_logic := '0';
    CZI29	: in std_logic := '0';
    CZI30	: in std_logic := '0';
    CZI31	: in std_logic := '0';
    CZI32	: in std_logic := '0';
    CZI33	: in std_logic := '0';
    CZI34	: in std_logic := '0';
    CZI35	: in std_logic := '0';
    CZI36	: in std_logic := '0';
    CZI37	: in std_logic := '0';
    CZI38	: in std_logic := '0';
    CZI39	: in std_logic := '0';
    CZI40	: in std_logic := '0';
    CZI41	: in std_logic := '0';
    CZI42	: in std_logic := '0';
    CZI43	: in std_logic := '0';
    CZI44	: in std_logic := '0';
    CZI45	: in std_logic := '0';
    CZI46	: in std_logic := '0';
    CZI47	: in std_logic := '0';
    CZI48	: in std_logic := '0';
    CZI49	: in std_logic := '0';
    CZI50	: in std_logic := '0';
    CZI51	: in std_logic := '0';
    CZI52	: in std_logic := '0';
    CZI53	: in std_logic := '0';
    CZI54	: in std_logic := '0';
    CZI55	: in std_logic := '0';
    CZI56	: in std_logic := '0';

    CZO1	: out std_logic := '0';
    CZO2	: out std_logic := '0';
    CZO3	: out std_logic := '0';
    CZO4	: out std_logic := '0';
    CZO5	: out std_logic := '0';
    CZO6	: out std_logic := '0';
    CZO7	: out std_logic := '0';
    CZO8	: out std_logic := '0';
    CZO9	: out std_logic := '0';
    CZO10	: out std_logic := '0';
    CZO11	: out std_logic := '0';
    CZO12	: out std_logic := '0';
    CZO13	: out std_logic := '0';
    CZO14	: out std_logic := '0';
    CZO15	: out std_logic := '0';
    CZO16	: out std_logic := '0';
    CZO17	: out std_logic := '0';
    CZO18	: out std_logic := '0';
    CZO19	: out std_logic := '0';
    CZO20	: out std_logic := '0';
    CZO21	: out std_logic := '0';
    CZO22	: out std_logic := '0';
    CZO23	: out std_logic := '0';
    CZO24	: out std_logic := '0';
    CZO25	: out std_logic := '0';
    CZO26	: out std_logic := '0';
    CZO27	: out std_logic := '0';
    CZO28	: out std_logic := '0';
    CZO29	: out std_logic := '0';
    CZO30	: out std_logic := '0';
    CZO31	: out std_logic := '0';
    CZO32	: out std_logic := '0';
    CZO33	: out std_logic := '0';
    CZO34	: out std_logic := '0';
    CZO35	: out std_logic := '0';
    CZO36	: out std_logic := '0';
    CZO37	: out std_logic := '0';
    CZO38	: out std_logic := '0';
    CZO39	: out std_logic := '0';
    CZO40	: out std_logic := '0';
    CZO41	: out std_logic := '0';
    CZO42	: out std_logic := '0';
    CZO43	: out std_logic := '0';
    CZO44	: out std_logic := '0';
    CZO45	: out std_logic := '0';
    CZO46	: out std_logic := '0';
    CZO47	: out std_logic := '0';
    CZO48	: out std_logic := '0';
    CZO49	: out std_logic := '0';
    CZO50	: out std_logic := '0';
    CZO51	: out std_logic := '0';
    CZO52	: out std_logic := '0';
    CZO53	: out std_logic := '0';
    CZO54	: out std_logic := '0';
    CZO55	: out std_logic := '0';
    CZO56	: out std_logic := '0';

    D1	: in std_logic := '0';
    D2	: in std_logic := '0';
    D3	: in std_logic := '0';
    D4	: in std_logic := '0';
    D5	: in std_logic := '0';
    D6	: in std_logic := '0';
    D7	: in std_logic := '0';
    D8	: in std_logic := '0';
    D9	: in std_logic := '0';
    D10	: in std_logic := '0';
    D11	: in std_logic := '0';
    D12	: in std_logic := '0';
    D13	: in std_logic := '0';
    D14	: in std_logic := '0';
    D15	: in std_logic := '0';
    D16	: in std_logic := '0';
    D17	: in std_logic := '0';
    D18	: in std_logic := '0';

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';

    Z1	: out std_logic := '0';
    Z2	: out std_logic := '0';
    Z3	: out std_logic := '0';
    Z4	: out std_logic := '0';
    Z5	: out std_logic := '0';
    Z6	: out std_logic := '0';
    Z7	: out std_logic := '0';
    Z8	: out std_logic := '0';
    Z9	: out std_logic := '0';
    Z10	: out std_logic := '0';
    Z11	: out std_logic := '0';
    Z12	: out std_logic := '0';
    Z13	: out std_logic := '0';
    Z14	: out std_logic := '0';
    Z15	: out std_logic := '0';
    Z16	: out std_logic := '0';
    Z17	: out std_logic := '0';
    Z18	: out std_logic := '0';
    Z19	: out std_logic := '0';
    Z20	: out std_logic := '0';
    Z21	: out std_logic := '0';
    Z22	: out std_logic := '0';
    Z23	: out std_logic := '0';
    Z24	: out std_logic := '0';
    Z25	: out std_logic := '0';
    Z26	: out std_logic := '0';
    Z27	: out std_logic := '0';
    Z28	: out std_logic := '0';
    Z29	: out std_logic := '0';
    Z30	: out std_logic := '0';
    Z31	: out std_logic := '0';
    Z32	: out std_logic := '0';
    Z33	: out std_logic := '0';
    Z34	: out std_logic := '0';
    Z35	: out std_logic := '0';
    Z36	: out std_logic := '0';
    Z37	: out std_logic := '0';
    Z38	: out std_logic := '0';
    Z39	: out std_logic := '0';
    Z40	: out std_logic := '0';
    Z41	: out std_logic := '0';
    Z42	: out std_logic := '0';
    Z43	: out std_logic := '0';
    Z44	: out std_logic := '0';
    Z45	: out std_logic := '0';
    Z46	: out std_logic := '0';
    Z47	: out std_logic := '0';
    Z48	: out std_logic := '0';
    Z49	: out std_logic := '0';
    Z50	: out std_logic := '0';
    Z51	: out std_logic := '0';
    Z52	: out std_logic := '0';
    Z53	: out std_logic := '0';
    Z54	: out std_logic := '0';
    Z55	: out std_logic := '0';
    Z56	: out std_logic := '0'
);
end component NX_DSP_L;

component NX_DSP_L_WRAP is
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A	: in std_logic_vector(23 downto 0) := (others => '0');
    B	: in std_logic_vector(17 downto 0) := (others => '0');
    C	: in std_logic_vector(35 downto 0) := (others => '0');

    CAI	: in std_logic_vector(23 downto 0) := (others => '0');
    CAO	: out std_logic_vector(23 downto 0) := (others => '0');
    CBI	: in std_logic_vector(17 downto 0) := (others => '0');
    CBO	: out std_logic_vector(17 downto 0) := (others => '0');

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO	: out std_logic := '0';
    CO37	: out std_logic := '0';
    CO57	: out std_logic := '0';

    CZI	: in std_logic_vector(55 downto 0) := (others => '0');
    CZO	: out std_logic_vector(55 downto 0) := (others => '0');

    D	: in std_logic_vector(17 downto 0) := (others => '0');

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0')
);
end component NX_DSP_L_WRAP;

component NX_DSP_L_SPLIT is
generic (
-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
------------------------------------------------------------------------- 
   SIGNED_MODE          : bit                    := '0';
   PRE_ADDER_OP         : bit                    := '0';       -- '0' = Additon, '1' = Subraction
   MUX_A                : bit                    := '0';       -- '0' = A input, '1' = CAI input
   MUX_B                : bit                    := '0';       -- '0' = B input, '1' = CBI input
   MUX_P                : bit                    := '0';       -- '0' for PRE_ADDER, '0' for B input
   MUX_X                : bit_vector(1 downto 0) := B"00";     -- Select X operand   "00" = C,
                                                               --                    "01" = CZI,
                                                               --                    "11" = SHFT(CZI) & C(11:0),
                                                               --                    "10" Select Z feedback
   MUX_Y                : bit                    := '0';       -- '0' Select MULT output, '1' for (B & A)
   MUX_CI               : bit                    := '0';       -- Select fabric input (not cascade)
   MUX_Z                : bit                    := '0';       -- Select ALU output
                                                               -- (not ALU input operand coming from PR_Y)

   Z_FEEDBACK_SHL12     : bit                    := '0';       -- '0' for No shift, '1' for 12-bit left shift
   ENABLE_SATURATION    : bit                    := '0';       -- '0' for Disable,  '1' for Enable
   SATURATION_RANK      : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB
                                                               --        on Z and CZO result
                                                               --(to define saturation and overflow)

   ALU_DYNAMIC_OP       : bit                    := '0';       -- '0' for Static,
                                                               -- '1' for Dynamic
                                                               -- (D6 ... D1 is not used for dynamic operation)
   CO_SEL               : bit                    := '0';       -- '0' for C0 = ALU(36), '1' for CO = ALU(48)

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
-------------------------------------------------------------------------
   PR_A_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on A input
   PR_A_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output
   PR_B_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on B input
   PR_B_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output

   PR_C_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_D_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_CI_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_P_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
   PR_X_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_Y_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

   PR_MULT_MUX             : bit                    := '0';   -- No pipe reg  -- Register inside MULT
   PR_ALU_MUX              : bit                    := '0';   -- No pipe reg  -- Register inside ALU
   PR_Z_MUX                : bit                    := '0';   -- Registered output

   PR_CO_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_OV_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
-------------------------------------------------------------------------
   ENABLE_PR_A_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_B_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_C_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_D_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CI_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_P_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_X_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Y_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_MULT_RST      : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_ALU_RST       : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Z_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CO_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_OV_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 

-------------------------------------------------------------------------
-- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
-------------------------------------------------------------------------
   ALU_OP                  : bit_vector(5 downto 0) := B"000000"; -- Addition = "000000", Subtract = "001010"
   ALU_MUX                 : bit                    := '0'        -- '0' for Don't swap ALU operands,
                                                                  -- '1' for ALU Swap operands
    );
port (
    CK	: IN std_logic := '0';
    R	: IN std_logic := '0';
    RZ	: IN std_logic := '0';
    WE	: IN std_logic := '0';

    CI	: IN std_logic := '0';
    A	: IN std_logic_vector(23 downto 0) := (others => '0');
    B	: IN std_logic_vector(17 downto 0) := (others => '0');
    C	: IN std_logic_vector(35 downto 0) := (others => '0');
    D	: IN std_logic_vector(17 downto 0) := (others => '0');
    CAI	: IN std_logic_vector(23 downto 0) := (others => '0');
    CBI	: IN std_logic_vector(17 downto 0) := (others => '0');
    CZI	: IN std_logic_vector(55 downto 0) := (others => '0');
    CCI	: IN std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0');
    CO	: OUT std_logic := '0';
    CO36	: OUT std_logic := '0';
    CO56	: OUT std_logic := '0';
    OVF	: OUT std_logic := '0';
    CAO	: OUT std_logic_vector(23 downto 0) := (others => '0');
    CBO	: OUT std_logic_vector(17 downto 0) := (others => '0');
    CZO	: OUT std_logic_vector(55 downto 0) := (others => '0');
    CCO	: OUT std_logic := '0'
  );
end component NX_DSP_L_SPLIT;

component NX_DSP is
generic (
    std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    A5	: in std_logic := '0';
    A6	: in std_logic := '0';
    A7	: in std_logic := '0';
    A8	: in std_logic := '0';
    A9	: in std_logic := '0';
    A10	: in std_logic := '0';
    A11	: in std_logic := '0';
    A12	: in std_logic := '0';
    A13	: in std_logic := '0';
    A14	: in std_logic := '0';
    A15	: in std_logic := '0';
    A16	: in std_logic := '0';
    A17	: in std_logic := '0';
    A18	: in std_logic := '0';
    A19	: in std_logic := '0';
    A20	: in std_logic := '0';
    A21	: in std_logic := '0';
    A22	: in std_logic := '0';
    A23	: in std_logic := '0';
    A24	: in std_logic := '0';

    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    B5	: in std_logic := '0';
    B6	: in std_logic := '0';
    B7	: in std_logic := '0';
    B8	: in std_logic := '0';
    B9	: in std_logic := '0';
    B10	: in std_logic := '0';
    B11	: in std_logic := '0';
    B12	: in std_logic := '0';
    B13	: in std_logic := '0';
    B14	: in std_logic := '0';
    B15	: in std_logic := '0';
    B16	: in std_logic := '0';
    B17	: in std_logic := '0';
    B18	: in std_logic := '0';

    C1	: in std_logic := '0';
    C2	: in std_logic := '0';
    C3	: in std_logic := '0';
    C4	: in std_logic := '0';
    C5	: in std_logic := '0';
    C6	: in std_logic := '0';
    C7	: in std_logic := '0';
    C8	: in std_logic := '0';
    C9	: in std_logic := '0';
    C10	: in std_logic := '0';
    C11	: in std_logic := '0';
    C12	: in std_logic := '0';
    C13	: in std_logic := '0';
    C14	: in std_logic := '0';
    C15	: in std_logic := '0';
    C16	: in std_logic := '0';
    C17	: in std_logic := '0';
    C18	: in std_logic := '0';
    C19	: in std_logic := '0';
    C20	: in std_logic := '0';
    C21	: in std_logic := '0';
    C22	: in std_logic := '0';
    C23	: in std_logic := '0';
    C24	: in std_logic := '0';
    C25	: in std_logic := '0';
    C26	: in std_logic := '0';
    C27	: in std_logic := '0';
    C28	: in std_logic := '0';
    C29	: in std_logic := '0';
    C30	: in std_logic := '0';
    C31	: in std_logic := '0';
    C32	: in std_logic := '0';
    C33	: in std_logic := '0';
    C34	: in std_logic := '0';
    C35	: in std_logic := '0';
    C36	: in std_logic := '0';

    CAI1	: in std_logic := '0';
    CAI2	: in std_logic := '0';
    CAI3	: in std_logic := '0';
    CAI4	: in std_logic := '0';
    CAI5	: in std_logic := '0';
    CAI6	: in std_logic := '0';
    CAI7	: in std_logic := '0';
    CAI8	: in std_logic := '0';
    CAI9	: in std_logic := '0';
    CAI10	: in std_logic := '0';
    CAI11	: in std_logic := '0';
    CAI12	: in std_logic := '0';
    CAI13	: in std_logic := '0';
    CAI14	: in std_logic := '0';
    CAI15	: in std_logic := '0';
    CAI16	: in std_logic := '0';
    CAI17	: in std_logic := '0';
    CAI18	: in std_logic := '0';

    CAO1	: out std_logic := '0';
    CAO2	: out std_logic := '0';
    CAO3	: out std_logic := '0';
    CAO4	: out std_logic := '0';
    CAO5	: out std_logic := '0';
    CAO6	: out std_logic := '0';
    CAO7	: out std_logic := '0';
    CAO8	: out std_logic := '0';
    CAO9	: out std_logic := '0';
    CAO10	: out std_logic := '0';
    CAO11	: out std_logic := '0';
    CAO12	: out std_logic := '0';
    CAO13	: out std_logic := '0';
    CAO14	: out std_logic := '0';
    CAO15	: out std_logic := '0';
    CAO16	: out std_logic := '0';
    CAO17	: out std_logic := '0';
    CAO18	: out std_logic := '0';

    CBI1	: in std_logic := '0';
    CBI2	: in std_logic := '0';
    CBI3	: in std_logic := '0';
    CBI4	: in std_logic := '0';
    CBI5	: in std_logic := '0';
    CBI6	: in std_logic := '0';
    CBI7	: in std_logic := '0';
    CBI8	: in std_logic := '0';
    CBI9	: in std_logic := '0';
    CBI10	: in std_logic := '0';
    CBI11	: in std_logic := '0';
    CBI12	: in std_logic := '0';
    CBI13	: in std_logic := '0';
    CBI14	: in std_logic := '0';
    CBI15	: in std_logic := '0';
    CBI16	: in std_logic := '0';
    CBI17	: in std_logic := '0';
    CBI18	: in std_logic := '0';

    CBO1	: out std_logic := '0';
    CBO2	: out std_logic := '0';
    CBO3	: out std_logic := '0';
    CBO4	: out std_logic := '0';
    CBO5	: out std_logic := '0';
    CBO6	: out std_logic := '0';
    CBO7	: out std_logic := '0';
    CBO8	: out std_logic := '0';
    CBO9	: out std_logic := '0';
    CBO10	: out std_logic := '0';
    CBO11	: out std_logic := '0';
    CBO12	: out std_logic := '0';
    CBO13	: out std_logic := '0';
    CBO14	: out std_logic := '0';
    CBO15	: out std_logic := '0';
    CBO16	: out std_logic := '0';
    CBO17	: out std_logic := '0';
    CBO18	: out std_logic := '0';

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO	: out std_logic := '0';
    CO37	: out std_logic := '0';
    CO49	: out std_logic := '0';

    CZI1	: in std_logic := '0';
    CZI2	: in std_logic := '0';
    CZI3	: in std_logic := '0';
    CZI4	: in std_logic := '0';
    CZI5	: in std_logic := '0';
    CZI6	: in std_logic := '0';
    CZI7	: in std_logic := '0';
    CZI8	: in std_logic := '0';
    CZI9	: in std_logic := '0';
    CZI10	: in std_logic := '0';
    CZI11	: in std_logic := '0';
    CZI12	: in std_logic := '0';
    CZI13	: in std_logic := '0';
    CZI14	: in std_logic := '0';
    CZI15	: in std_logic := '0';
    CZI16	: in std_logic := '0';
    CZI17	: in std_logic := '0';
    CZI18	: in std_logic := '0';
    CZI19	: in std_logic := '0';
    CZI20	: in std_logic := '0';
    CZI21	: in std_logic := '0';
    CZI22	: in std_logic := '0';
    CZI23	: in std_logic := '0';
    CZI24	: in std_logic := '0';
    CZI25	: in std_logic := '0';
    CZI26	: in std_logic := '0';
    CZI27	: in std_logic := '0';
    CZI28	: in std_logic := '0';
    CZI29	: in std_logic := '0';
    CZI30	: in std_logic := '0';
    CZI31	: in std_logic := '0';
    CZI32	: in std_logic := '0';
    CZI33	: in std_logic := '0';
    CZI34	: in std_logic := '0';
    CZI35	: in std_logic := '0';
    CZI36	: in std_logic := '0';
    CZI37	: in std_logic := '0';
    CZI38	: in std_logic := '0';
    CZI39	: in std_logic := '0';
    CZI40	: in std_logic := '0';
    CZI41	: in std_logic := '0';
    CZI42	: in std_logic := '0';
    CZI43	: in std_logic := '0';
    CZI44	: in std_logic := '0';
    CZI45	: in std_logic := '0';
    CZI46	: in std_logic := '0';
    CZI47	: in std_logic := '0';
    CZI48	: in std_logic := '0';
    CZI49	: in std_logic := '0';
    CZI50	: in std_logic := '0';
    CZI51	: in std_logic := '0';
    CZI52	: in std_logic := '0';
    CZI53	: in std_logic := '0';
    CZI54	: in std_logic := '0';
    CZI55	: in std_logic := '0';
    CZI56	: in std_logic := '0';

    CZO1	: out std_logic := '0';
    CZO2	: out std_logic := '0';
    CZO3	: out std_logic := '0';
    CZO4	: out std_logic := '0';
    CZO5	: out std_logic := '0';
    CZO6	: out std_logic := '0';
    CZO7	: out std_logic := '0';
    CZO8	: out std_logic := '0';
    CZO9	: out std_logic := '0';
    CZO10	: out std_logic := '0';
    CZO11	: out std_logic := '0';
    CZO12	: out std_logic := '0';
    CZO13	: out std_logic := '0';
    CZO14	: out std_logic := '0';
    CZO15	: out std_logic := '0';
    CZO16	: out std_logic := '0';
    CZO17	: out std_logic := '0';
    CZO18	: out std_logic := '0';
    CZO19	: out std_logic := '0';
    CZO20	: out std_logic := '0';
    CZO21	: out std_logic := '0';
    CZO22	: out std_logic := '0';
    CZO23	: out std_logic := '0';
    CZO24	: out std_logic := '0';
    CZO25	: out std_logic := '0';
    CZO26	: out std_logic := '0';
    CZO27	: out std_logic := '0';
    CZO28	: out std_logic := '0';
    CZO29	: out std_logic := '0';
    CZO30	: out std_logic := '0';
    CZO31	: out std_logic := '0';
    CZO32	: out std_logic := '0';
    CZO33	: out std_logic := '0';
    CZO34	: out std_logic := '0';
    CZO35	: out std_logic := '0';
    CZO36	: out std_logic := '0';
    CZO37	: out std_logic := '0';
    CZO38	: out std_logic := '0';
    CZO39	: out std_logic := '0';
    CZO40	: out std_logic := '0';
    CZO41	: out std_logic := '0';
    CZO42	: out std_logic := '0';
    CZO43	: out std_logic := '0';
    CZO44	: out std_logic := '0';
    CZO45	: out std_logic := '0';
    CZO46	: out std_logic := '0';
    CZO47	: out std_logic := '0';
    CZO48	: out std_logic := '0';
    CZO49	: out std_logic := '0';
    CZO50	: out std_logic := '0';
    CZO51	: out std_logic := '0';
    CZO52	: out std_logic := '0';
    CZO53	: out std_logic := '0';
    CZO54	: out std_logic := '0';
    CZO55	: out std_logic := '0';
    CZO56	: out std_logic := '0';

    D1	: in std_logic := '0';
    D2	: in std_logic := '0';
    D3	: in std_logic := '0';
    D4	: in std_logic := '0';
    D5	: in std_logic := '0';
    D6	: in std_logic := '0';
    D7	: in std_logic := '0';
    D8	: in std_logic := '0';
    D9	: in std_logic := '0';
    D10	: in std_logic := '0';
    D11	: in std_logic := '0';
    D12	: in std_logic := '0';
    D13	: in std_logic := '0';
    D14	: in std_logic := '0';
    D15	: in std_logic := '0';
    D16	: in std_logic := '0';
    D17	: in std_logic := '0';
    D18	: in std_logic := '0';

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';

    Z1	: out std_logic := '0';
    Z2	: out std_logic := '0';
    Z3	: out std_logic := '0';
    Z4	: out std_logic := '0';
    Z5	: out std_logic := '0';
    Z6	: out std_logic := '0';
    Z7	: out std_logic := '0';
    Z8	: out std_logic := '0';
    Z9	: out std_logic := '0';
    Z10	: out std_logic := '0';
    Z11	: out std_logic := '0';
    Z12	: out std_logic := '0';
    Z13	: out std_logic := '0';
    Z14	: out std_logic := '0';
    Z15	: out std_logic := '0';
    Z16	: out std_logic := '0';
    Z17	: out std_logic := '0';
    Z18	: out std_logic := '0';
    Z19	: out std_logic := '0';
    Z20	: out std_logic := '0';
    Z21	: out std_logic := '0';
    Z22	: out std_logic := '0';
    Z23	: out std_logic := '0';
    Z24	: out std_logic := '0';
    Z25	: out std_logic := '0';
    Z26	: out std_logic := '0';
    Z27	: out std_logic := '0';
    Z28	: out std_logic := '0';
    Z29	: out std_logic := '0';
    Z30	: out std_logic := '0';
    Z31	: out std_logic := '0';
    Z32	: out std_logic := '0';
    Z33	: out std_logic := '0';
    Z34	: out std_logic := '0';
    Z35	: out std_logic := '0';
    Z36	: out std_logic := '0';
    Z37	: out std_logic := '0';
    Z38	: out std_logic := '0';
    Z39	: out std_logic := '0';
    Z40	: out std_logic := '0';
    Z41	: out std_logic := '0';
    Z42	: out std_logic := '0';
    Z43	: out std_logic := '0';
    Z44	: out std_logic := '0';
    Z45	: out std_logic := '0';
    Z46	: out std_logic := '0';
    Z47	: out std_logic := '0';
    Z48	: out std_logic := '0';
    Z49	: out std_logic := '0';
    Z50	: out std_logic := '0';
    Z51	: out std_logic := '0';
    Z52	: out std_logic := '0';
    Z53	: out std_logic := '0';
    Z54	: out std_logic := '0';
    Z55	: out std_logic := '0';
    Z56	: out std_logic := '0'
);
end component NX_DSP;

component NX_DSP_WRAP is
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A	: in std_logic_vector(23 downto 0) := (others => '0');
    B	: in std_logic_vector(17 downto 0) := (others => '0');
    C	: in std_logic_vector(35 downto 0) := (others => '0');

    CAI	: in std_logic_vector(17 downto 0) := (others => '0');
    CAO	: out std_logic_vector(17 downto 0) := (others => '0');
    CBI	: in std_logic_vector(17 downto 0) := (others => '0');
    CBO	: out std_logic_vector(17 downto 0) := (others => '0');

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO	: out std_logic := '0';
    CO37	: out std_logic := '0';
    CO49	: out std_logic := '0';

    CZI	: in std_logic_vector(55 downto 0) := (others => '0');
    CZO	: out std_logic_vector(55 downto 0) := (others => '0');

    D	: in std_logic_vector(17 downto 0) := (others => '0');

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0')
);
end component NX_DSP_WRAP;

component NX_DSP_SPLIT is
generic (
-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
------------------------------------------------------------------------- 
   SIGNED_MODE          : bit                    := '0';
   PRE_ADDER_OP         : bit                    := '0';       -- '0' = Additon, '1' = Subraction
   MUX_A                : bit                    := '0';       -- '0' = A input, '1' = CAI input
   MUX_B                : bit                    := '0';       -- '0' = B input, '1' = CBI input
   MUX_P                : bit                    := '0';       -- '0' for PRE_ADDER, '0' for B input
   MUX_X                : bit_vector(1 downto 0) := B"00";     -- Select X operand   "00" = C,
                                                               --                    "01" = CZI,
                                                               --                    "11" = SHFT(CZI) & C(11:0),
                                                               --                    "10" Select Z feedback
   MUX_Y                : bit                    := '0';       -- '0' Select MULT output, '1' for (B & A)
   MUX_CI               : bit                    := '0';       -- Select fabric input (not cascade)
   MUX_Z                : bit                    := '0';       -- Select ALU output
                                                               -- (not ALU input operand coming from PR_Y)

   Z_FEEDBACK_SHL12     : bit                    := '0';       -- '0' for No shift, '1' for 12-bit left shift
   ENABLE_SATURATION    : bit                    := '0';       -- '0' for Disable,  '1' for Enable
   SATURATION_RANK      : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB
                                                               --        on Z and CZO result
                                                               --(to define saturation and overflow)

   ALU_DYNAMIC_OP       : bit                    := '0';       -- '0' for Static,
                                                               -- '1' for Dynamic
                                                               -- (D6 ... D1 is not used for dynamic operation)
   CO_SEL               : bit                    := '0';       -- '0' for C0 = ALU(36), '1' for CO = ALU(48)

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
-------------------------------------------------------------------------
   PR_A_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on A input
   PR_A_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output
   PR_B_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on B input
   PR_B_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output

   PR_C_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_D_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_CI_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_P_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
   PR_X_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_Y_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

   PR_MULT_MUX             : bit                    := '0';   -- No pipe reg  -- Register inside MULT
   PR_ALU_MUX              : bit                    := '0';   -- No pipe reg  -- Register inside ALU
   PR_Z_MUX                : bit                    := '0';   -- Registered output

   PR_CO_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_OV_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
-------------------------------------------------------------------------
   ENABLE_PR_A_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_B_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_C_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_D_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CI_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_P_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_X_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Y_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_MULT_RST      : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_ALU_RST       : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Z_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CO_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_OV_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 

-------------------------------------------------------------------------
-- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
-------------------------------------------------------------------------
   ALU_OP                  : bit_vector(5 downto 0) := B"000000"; -- Addition = "000000", Subtract = "001010"
   ALU_MUX                 : bit                    := '0'        -- '0' for Don't swap ALU operands,
                                                                  -- '1' for ALU Swap operands
    );
port (
    CK	: IN std_logic := '0';
    R	: IN std_logic := '0';
    RZ	: IN std_logic := '0';
    WE	: IN std_logic := '0';

    CI	: IN std_logic := '0';
    A	: IN std_logic_vector(23 downto 0) := (others => '0');
    B	: IN std_logic_vector(17 downto 0) := (others => '0');
    C	: IN std_logic_vector(35 downto 0) := (others => '0');
    D	: IN std_logic_vector(17 downto 0) := (others => '0');
    CAI	: IN std_logic_vector(17 downto 0) := (others => '0');
    CBI	: IN std_logic_vector(17 downto 0) := (others => '0');
    CZI	: IN std_logic_vector(55 downto 0) := (others => '0');
    CCI	: IN std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0');
    CO	: OUT std_logic := '0';
    CO36	: OUT std_logic := '0';
    CO48	: OUT std_logic := '0';
    OVF	: OUT std_logic := '0';
    CAO	: OUT std_logic_vector(17 downto 0) := (others => '0');
    CBO	: OUT std_logic_vector(17 downto 0) := (others => '0');
    CZO	: OUT std_logic_vector(55 downto 0) := (others => '0');
    CCO	: OUT std_logic := '0'
  );
end component NX_DSP_SPLIT;

component NX_DSPDPRAM_FULL_U is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    dsp0_clk_i	: in std_logic := '0';
    dsp0_rst_i	: in std_logic := '0';
    dsp0_rstz_i	: in std_logic := '0';
    dsp0_we_i	: in std_logic := '0';
    dsp0_wez_i	: in std_logic := '0';
    dsp0_cy_i	: in std_logic := '0';
    dsp0_a_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dsp0_b_i	: in std_logic_vector(17 downto 0) := (others => '0');
    dsp0_c_i	: in std_logic_vector(35 downto 0) := (others => '0');
    dsp0_d_i	: in std_logic_vector(17 downto 0) := (others => '0');

    dsp0_z_o	: out std_logic_vector(55 downto 0) := (others => '0');
    dsp0_cy_o	: out std_logic := '0';
    dsp0_cy42_o	: out std_logic := '0';
    dsp0_cy56_o	: out std_logic := '0';
    dsp0_ovf_o	: out std_logic := '0';

    dsp1_clk_i	: in std_logic := '0';
    dsp1_rst_i	: in std_logic := '0';
    dsp1_rstz_i	: in std_logic := '0';
    dsp1_we_i	: in std_logic := '0';
    dsp1_wez_i	: in std_logic := '0';
    dsp1_cy_i	: in std_logic := '0';
    dsp1_a_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dsp1_b_i	: in std_logic_vector(17 downto 0) := (others => '0');
    dsp1_c_i	: in std_logic_vector(35 downto 0) := (others => '0');
    dsp1_d_i	: in std_logic_vector(17 downto 0) := (others => '0');

    dsp1_z_o	: out std_logic_vector(55 downto 0) := (others => '0');
    dsp1_cy_o	: out std_logic := '0';
    dsp1_cy42_o	: out std_logic := '0';
    dsp1_cy56_o	: out std_logic := '0';
    dsp1_ovf_o	: out std_logic := '0';

    dpram_clkmem0_i	: in std_logic := '0';
    dpram_rst0_i	: in std_logic := '0';
    dpram_cs0_i	: in std_logic := '0';
    dpram_we0_i	: in std_logic := '0';
    dpram_addr0_i	: in std_logic_vector(15 downto 0) := (others => '0');
    dpram_din0_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dpram_dout0_o	: out std_logic_vector(23 downto 0) := (others => '0');
    dpram_ecc_corrected0_o	: out std_logic := '0';
    dpram_ecc_uncorrected0_o	: out std_logic := '0';

    dpram_clkmem1_i	: in std_logic := '0';
    dpram_rst1_i	: in std_logic := '0';
    dpram_cs1_i	: in std_logic := '0';
    dpram_we1_i	: in std_logic := '0';
    dpram_addr1_i	: in std_logic_vector(15 downto 0) := (others => '0');
    dpram_din1_i	: in std_logic_vector(23 downto 0) := (others => '0');
    dpram_dout1_o	: out std_logic_vector(23 downto 0) := (others => '0');
    dpram_ecc_corrected1_o	: out std_logic := '0';
    dpram_ecc_uncorrected1_o	: out std_logic := '0'
);
end component NX_DSPDPRAM_FULL_U;

component NX_DSP_U_BOX is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    A5	: in std_logic := '0';
    A6	: in std_logic := '0';
    A7	: in std_logic := '0';
    A8	: in std_logic := '0';
    A9	: in std_logic := '0';
    A10	: in std_logic := '0';
    A11	: in std_logic := '0';
    A12	: in std_logic := '0';
    A13	: in std_logic := '0';
    A14	: in std_logic := '0';
    A15	: in std_logic := '0';
    A16	: in std_logic := '0';
    A17	: in std_logic := '0';
    A18	: in std_logic := '0';
    A19	: in std_logic := '0';
    A20	: in std_logic := '0';
    A21	: in std_logic := '0';
    A22	: in std_logic := '0';
    A23	: in std_logic := '0';
    A24	: in std_logic := '0';

    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    B5	: in std_logic := '0';
    B6	: in std_logic := '0';
    B7	: in std_logic := '0';
    B8	: in std_logic := '0';
    B9	: in std_logic := '0';
    B10	: in std_logic := '0';
    B11	: in std_logic := '0';
    B12	: in std_logic := '0';
    B13	: in std_logic := '0';
    B14	: in std_logic := '0';
    B15	: in std_logic := '0';
    B16	: in std_logic := '0';
    B17	: in std_logic := '0';
    B18	: in std_logic := '0';

    C1	: in std_logic := '0';
    C2	: in std_logic := '0';
    C3	: in std_logic := '0';
    C4	: in std_logic := '0';
    C5	: in std_logic := '0';
    C6	: in std_logic := '0';
    C7	: in std_logic := '0';
    C8	: in std_logic := '0';
    C9	: in std_logic := '0';
    C10	: in std_logic := '0';
    C11	: in std_logic := '0';
    C12	: in std_logic := '0';
    C13	: in std_logic := '0';
    C14	: in std_logic := '0';
    C15	: in std_logic := '0';
    C16	: in std_logic := '0';
    C17	: in std_logic := '0';
    C18	: in std_logic := '0';
    C19	: in std_logic := '0';
    C20	: in std_logic := '0';
    C21	: in std_logic := '0';
    C22	: in std_logic := '0';
    C23	: in std_logic := '0';
    C24	: in std_logic := '0';
    C25	: in std_logic := '0';
    C26	: in std_logic := '0';
    C27	: in std_logic := '0';
    C28	: in std_logic := '0';
    C29	: in std_logic := '0';
    C30	: in std_logic := '0';
    C31	: in std_logic := '0';
    C32	: in std_logic := '0';
    C33	: in std_logic := '0';
    C34	: in std_logic := '0';
    C35	: in std_logic := '0';
    C36	: in std_logic := '0';

    CAI1	: in std_logic := '0';
    CAI2	: in std_logic := '0';
    CAI3	: in std_logic := '0';
    CAI4	: in std_logic := '0';
    CAI5	: in std_logic := '0';
    CAI6	: in std_logic := '0';
    CAI7	: in std_logic := '0';
    CAI8	: in std_logic := '0';
    CAI9	: in std_logic := '0';
    CAI10	: in std_logic := '0';
    CAI11	: in std_logic := '0';
    CAI12	: in std_logic := '0';
    CAI13	: in std_logic := '0';
    CAI14	: in std_logic := '0';
    CAI15	: in std_logic := '0';
    CAI16	: in std_logic := '0';
    CAI17	: in std_logic := '0';
    CAI18	: in std_logic := '0';
    CAI19	: in std_logic := '0';
    CAI20	: in std_logic := '0';
    CAI21	: in std_logic := '0';
    CAI22	: in std_logic := '0';
    CAI23	: in std_logic := '0';
    CAI24	: in std_logic := '0';

    CAO1	: out std_logic := '0';
    CAO2	: out std_logic := '0';
    CAO3	: out std_logic := '0';
    CAO4	: out std_logic := '0';
    CAO5	: out std_logic := '0';
    CAO6	: out std_logic := '0';
    CAO7	: out std_logic := '0';
    CAO8	: out std_logic := '0';
    CAO9	: out std_logic := '0';
    CAO10	: out std_logic := '0';
    CAO11	: out std_logic := '0';
    CAO12	: out std_logic := '0';
    CAO13	: out std_logic := '0';
    CAO14	: out std_logic := '0';
    CAO15	: out std_logic := '0';
    CAO16	: out std_logic := '0';
    CAO17	: out std_logic := '0';
    CAO18	: out std_logic := '0';
    CAO19	: out std_logic := '0';
    CAO20	: out std_logic := '0';
    CAO21	: out std_logic := '0';
    CAO22	: out std_logic := '0';
    CAO23	: out std_logic := '0';
    CAO24	: out std_logic := '0';

    CBI1	: in std_logic := '0';
    CBI2	: in std_logic := '0';
    CBI3	: in std_logic := '0';
    CBI4	: in std_logic := '0';
    CBI5	: in std_logic := '0';
    CBI6	: in std_logic := '0';
    CBI7	: in std_logic := '0';
    CBI8	: in std_logic := '0';
    CBI9	: in std_logic := '0';
    CBI10	: in std_logic := '0';
    CBI11	: in std_logic := '0';
    CBI12	: in std_logic := '0';
    CBI13	: in std_logic := '0';
    CBI14	: in std_logic := '0';
    CBI15	: in std_logic := '0';
    CBI16	: in std_logic := '0';
    CBI17	: in std_logic := '0';
    CBI18	: in std_logic := '0';

    CBO1	: out std_logic := '0';
    CBO2	: out std_logic := '0';
    CBO3	: out std_logic := '0';
    CBO4	: out std_logic := '0';
    CBO5	: out std_logic := '0';
    CBO6	: out std_logic := '0';
    CBO7	: out std_logic := '0';
    CBO8	: out std_logic := '0';
    CBO9	: out std_logic := '0';
    CBO10	: out std_logic := '0';
    CBO11	: out std_logic := '0';
    CBO12	: out std_logic := '0';
    CBO13	: out std_logic := '0';
    CBO14	: out std_logic := '0';
    CBO15	: out std_logic := '0';
    CBO16	: out std_logic := '0';
    CBO17	: out std_logic := '0';
    CBO18	: out std_logic := '0';

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    RESERVED: out std_logic;
    CO43	: out std_logic := '0';
    CO57	: out std_logic := '0';

    CZI1	: in std_logic := '0';
    CZI2	: in std_logic := '0';
    CZI3	: in std_logic := '0';
    CZI4	: in std_logic := '0';
    CZI5	: in std_logic := '0';
    CZI6	: in std_logic := '0';
    CZI7	: in std_logic := '0';
    CZI8	: in std_logic := '0';
    CZI9	: in std_logic := '0';
    CZI10	: in std_logic := '0';
    CZI11	: in std_logic := '0';
    CZI12	: in std_logic := '0';
    CZI13	: in std_logic := '0';
    CZI14	: in std_logic := '0';
    CZI15	: in std_logic := '0';
    CZI16	: in std_logic := '0';
    CZI17	: in std_logic := '0';
    CZI18	: in std_logic := '0';
    CZI19	: in std_logic := '0';
    CZI20	: in std_logic := '0';
    CZI21	: in std_logic := '0';
    CZI22	: in std_logic := '0';
    CZI23	: in std_logic := '0';
    CZI24	: in std_logic := '0';
    CZI25	: in std_logic := '0';
    CZI26	: in std_logic := '0';
    CZI27	: in std_logic := '0';
    CZI28	: in std_logic := '0';
    CZI29	: in std_logic := '0';
    CZI30	: in std_logic := '0';
    CZI31	: in std_logic := '0';
    CZI32	: in std_logic := '0';
    CZI33	: in std_logic := '0';
    CZI34	: in std_logic := '0';
    CZI35	: in std_logic := '0';
    CZI36	: in std_logic := '0';
    CZI37	: in std_logic := '0';
    CZI38	: in std_logic := '0';
    CZI39	: in std_logic := '0';
    CZI40	: in std_logic := '0';
    CZI41	: in std_logic := '0';
    CZI42	: in std_logic := '0';
    CZI43	: in std_logic := '0';
    CZI44	: in std_logic := '0';
    CZI45	: in std_logic := '0';
    CZI46	: in std_logic := '0';
    CZI47	: in std_logic := '0';
    CZI48	: in std_logic := '0';
    CZI49	: in std_logic := '0';
    CZI50	: in std_logic := '0';
    CZI51	: in std_logic := '0';
    CZI52	: in std_logic := '0';
    CZI53	: in std_logic := '0';
    CZI54	: in std_logic := '0';
    CZI55	: in std_logic := '0';
    CZI56	: in std_logic := '0';

    CZO1	: out std_logic := '0';
    CZO2	: out std_logic := '0';
    CZO3	: out std_logic := '0';
    CZO4	: out std_logic := '0';
    CZO5	: out std_logic := '0';
    CZO6	: out std_logic := '0';
    CZO7	: out std_logic := '0';
    CZO8	: out std_logic := '0';
    CZO9	: out std_logic := '0';
    CZO10	: out std_logic := '0';
    CZO11	: out std_logic := '0';
    CZO12	: out std_logic := '0';
    CZO13	: out std_logic := '0';
    CZO14	: out std_logic := '0';
    CZO15	: out std_logic := '0';
    CZO16	: out std_logic := '0';
    CZO17	: out std_logic := '0';
    CZO18	: out std_logic := '0';
    CZO19	: out std_logic := '0';
    CZO20	: out std_logic := '0';
    CZO21	: out std_logic := '0';
    CZO22	: out std_logic := '0';
    CZO23	: out std_logic := '0';
    CZO24	: out std_logic := '0';
    CZO25	: out std_logic := '0';
    CZO26	: out std_logic := '0';
    CZO27	: out std_logic := '0';
    CZO28	: out std_logic := '0';
    CZO29	: out std_logic := '0';
    CZO30	: out std_logic := '0';
    CZO31	: out std_logic := '0';
    CZO32	: out std_logic := '0';
    CZO33	: out std_logic := '0';
    CZO34	: out std_logic := '0';
    CZO35	: out std_logic := '0';
    CZO36	: out std_logic := '0';
    CZO37	: out std_logic := '0';
    CZO38	: out std_logic := '0';
    CZO39	: out std_logic := '0';
    CZO40	: out std_logic := '0';
    CZO41	: out std_logic := '0';
    CZO42	: out std_logic := '0';
    CZO43	: out std_logic := '0';
    CZO44	: out std_logic := '0';
    CZO45	: out std_logic := '0';
    CZO46	: out std_logic := '0';
    CZO47	: out std_logic := '0';
    CZO48	: out std_logic := '0';
    CZO49	: out std_logic := '0';
    CZO50	: out std_logic := '0';
    CZO51	: out std_logic := '0';
    CZO52	: out std_logic := '0';
    CZO53	: out std_logic := '0';
    CZO54	: out std_logic := '0';
    CZO55	: out std_logic := '0';
    CZO56	: out std_logic := '0';

    D1	: in std_logic := '0';
    D2	: in std_logic := '0';
    D3	: in std_logic := '0';
    D4	: in std_logic := '0';
    D5	: in std_logic := '0';
    D6	: in std_logic := '0';
    D7	: in std_logic := '0';
    D8	: in std_logic := '0';
    D9	: in std_logic := '0';
    D10	: in std_logic := '0';
    D11	: in std_logic := '0';
    D12	: in std_logic := '0';
    D13	: in std_logic := '0';
    D14	: in std_logic := '0';
    D15	: in std_logic := '0';
    D16	: in std_logic := '0';
    D17	: in std_logic := '0';
    D18	: in std_logic := '0';

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEZ	: in std_logic := '0';

    Z1	: out std_logic := '0';
    Z2	: out std_logic := '0';
    Z3	: out std_logic := '0';
    Z4	: out std_logic := '0';
    Z5	: out std_logic := '0';
    Z6	: out std_logic := '0';
    Z7	: out std_logic := '0';
    Z8	: out std_logic := '0';
    Z9	: out std_logic := '0';
    Z10	: out std_logic := '0';
    Z11	: out std_logic := '0';
    Z12	: out std_logic := '0';
    Z13	: out std_logic := '0';
    Z14	: out std_logic := '0';
    Z15	: out std_logic := '0';
    Z16	: out std_logic := '0';
    Z17	: out std_logic := '0';
    Z18	: out std_logic := '0';
    Z19	: out std_logic := '0';
    Z20	: out std_logic := '0';
    Z21	: out std_logic := '0';
    Z22	: out std_logic := '0';
    Z23	: out std_logic := '0';
    Z24	: out std_logic := '0';
    Z25	: out std_logic := '0';
    Z26	: out std_logic := '0';
    Z27	: out std_logic := '0';
    Z28	: out std_logic := '0';
    Z29	: out std_logic := '0';
    Z30	: out std_logic := '0';
    Z31	: out std_logic := '0';
    Z32	: out std_logic := '0';
    Z33	: out std_logic := '0';
    Z34	: out std_logic := '0';
    Z35	: out std_logic := '0';
    Z36	: out std_logic := '0';
    Z37	: out std_logic := '0';
    Z38	: out std_logic := '0';
    Z39	: out std_logic := '0';
    Z40	: out std_logic := '0';
    Z41	: out std_logic := '0';
    Z42	: out std_logic := '0';
    Z43	: out std_logic := '0';
    Z44	: out std_logic := '0';
    Z45	: out std_logic := '0';
    Z46	: out std_logic := '0';
    Z47	: out std_logic := '0';
    Z48	: out std_logic := '0';
    Z49	: out std_logic := '0';
    Z50	: out std_logic := '0';
    Z51	: out std_logic := '0';
    Z52	: out std_logic := '0';
    Z53	: out std_logic := '0';
    Z54	: out std_logic := '0';
    Z55	: out std_logic := '0';
    Z56	: out std_logic := '0'
);
end component NX_DSP_U_BOX;

component NX_RAM_U_BOX is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    ACK	: in std_logic := '0';
    BCK	: in std_logic := '0';

    AI1	: in std_logic := '0';
    AI2	: in std_logic := '0';
    AI3	: in std_logic := '0';
    AI4	: in std_logic := '0';
    AI5	: in std_logic := '0';
    AI6	: in std_logic := '0';
    AI7	: in std_logic := '0';
    AI8	: in std_logic := '0';
    AI9	: in std_logic := '0';
    AI10	: in std_logic := '0';
    AI11	: in std_logic := '0';
    AI12	: in std_logic := '0';
    AI13	: in std_logic := '0';
    AI14	: in std_logic := '0';
    AI15	: in std_logic := '0';
    AI16	: in std_logic := '0';
    AI17	: in std_logic := '0';
    AI18	: in std_logic := '0';
    AI19	: in std_logic := '0';
    AI20	: in std_logic := '0';
    AI21	: in std_logic := '0';
    AI22	: in std_logic := '0';
    AI23	: in std_logic := '0';
    AI24	: in std_logic := '0';

    BI1	: in std_logic := '0';
    BI2	: in std_logic := '0';
    BI3	: in std_logic := '0';
    BI4	: in std_logic := '0';
    BI5	: in std_logic := '0';
    BI6	: in std_logic := '0';
    BI7	: in std_logic := '0';
    BI8	: in std_logic := '0';
    BI9	: in std_logic := '0';
    BI10	: in std_logic := '0';
    BI11	: in std_logic := '0';
    BI12	: in std_logic := '0';
    BI13	: in std_logic := '0';
    BI14	: in std_logic := '0';
    BI15	: in std_logic := '0';
    BI16	: in std_logic := '0';
    BI17	: in std_logic := '0';
    BI18	: in std_logic := '0';
    BI19	: in std_logic := '0';
    BI20	: in std_logic := '0';
    BI21	: in std_logic := '0';
    BI22	: in std_logic := '0';
    BI23	: in std_logic := '0';
    BI24	: in std_logic := '0';

    ACOR	: out std_logic := '0';
    AERR	: out std_logic := '0';
    BCOR	: out std_logic := '0';
    BERR	: out std_logic := '0';

    AO1	: out std_logic := '0';
    AO2	: out std_logic := '0';
    AO3	: out std_logic := '0';
    AO4	: out std_logic := '0';
    AO5	: out std_logic := '0';
    AO6	: out std_logic := '0';
    AO7	: out std_logic := '0';
    AO8	: out std_logic := '0';
    AO9	: out std_logic := '0';
    AO10	: out std_logic := '0';
    AO11	: out std_logic := '0';
    AO12	: out std_logic := '0';
    AO13	: out std_logic := '0';
    AO14	: out std_logic := '0';
    AO15	: out std_logic := '0';
    AO16	: out std_logic := '0';
    AO17	: out std_logic := '0';
    AO18	: out std_logic := '0';
    AO19	: out std_logic := '0';
    AO20	: out std_logic := '0';
    AO21	: out std_logic := '0';
    AO22	: out std_logic := '0';
    AO23	: out std_logic := '0';
    AO24	: out std_logic := '0';

    BO1	: out std_logic := '0';
    BO2	: out std_logic := '0';
    BO3	: out std_logic := '0';
    BO4	: out std_logic := '0';
    BO5	: out std_logic := '0';
    BO6	: out std_logic := '0';
    BO7	: out std_logic := '0';
    BO8	: out std_logic := '0';
    BO9	: out std_logic := '0';
    BO10	: out std_logic := '0';
    BO11	: out std_logic := '0';
    BO12	: out std_logic := '0';
    BO13	: out std_logic := '0';
    BO14	: out std_logic := '0';
    BO15	: out std_logic := '0';
    BO16	: out std_logic := '0';
    BO17	: out std_logic := '0';
    BO18	: out std_logic := '0';
    BO19	: out std_logic := '0';
    BO20	: out std_logic := '0';
    BO21	: out std_logic := '0';
    BO22	: out std_logic := '0';
    BO23	: out std_logic := '0';
    BO24	: out std_logic := '0';

    AA1	: in std_logic := '0';
    AA2	: in std_logic := '0';
    AA3	: in std_logic := '0';
    AA4	: in std_logic := '0';
    AA5	: in std_logic := '0';
    AA6	: in std_logic := '0';
    AA7	: in std_logic := '0';
    AA8	: in std_logic := '0';
    AA9	: in std_logic := '0';
    AA10	: in std_logic := '0';
    AA11	: in std_logic := '0';
    AA12	: in std_logic := '0';
    AA13	: in std_logic := '0';
    AA14	: in std_logic := '0';
    AA15	: in std_logic := '0';
    AA16	: in std_logic := '0';

    ACS	: in std_logic := '0';
    AWE	: in std_logic := '0';
    AR	: in std_logic := '0';

    BA1	: in std_logic := '0';
    BA2	: in std_logic := '0';
    BA3	: in std_logic := '0';
    BA4	: in std_logic := '0';
    BA5	: in std_logic := '0';
    BA6	: in std_logic := '0';
    BA7	: in std_logic := '0';
    BA8	: in std_logic := '0';
    BA9	: in std_logic := '0';
    BA10	: in std_logic := '0';
    BA11	: in std_logic := '0';
    BA12	: in std_logic := '0';
    BA13	: in std_logic := '0';
    BA14	: in std_logic := '0';
    BA15	: in std_logic := '0';
    BA16	: in std_logic := '0';

    BCS	: in std_logic := '0';
    BWE	: in std_logic := '0';
    BR	: in std_logic := '0'
);
end component NX_RAM_U_BOX;

component NX_DSP_U is
generic (
        std_mode    : string                  := "";                             -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
        raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
        raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
        raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
        raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
    );
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    A5	: in std_logic := '0';
    A6	: in std_logic := '0';
    A7	: in std_logic := '0';
    A8	: in std_logic := '0';
    A9	: in std_logic := '0';
    A10	: in std_logic := '0';
    A11	: in std_logic := '0';
    A12	: in std_logic := '0';
    A13	: in std_logic := '0';
    A14	: in std_logic := '0';
    A15	: in std_logic := '0';
    A16	: in std_logic := '0';
    A17	: in std_logic := '0';
    A18	: in std_logic := '0';
    A19	: in std_logic := '0';
    A20	: in std_logic := '0';
    A21	: in std_logic := '0';
    A22	: in std_logic := '0';
    A23	: in std_logic := '0';
    A24	: in std_logic := '0';

    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    B5	: in std_logic := '0';
    B6	: in std_logic := '0';
    B7	: in std_logic := '0';
    B8	: in std_logic := '0';
    B9	: in std_logic := '0';
    B10	: in std_logic := '0';
    B11	: in std_logic := '0';
    B12	: in std_logic := '0';
    B13	: in std_logic := '0';
    B14	: in std_logic := '0';
    B15	: in std_logic := '0';
    B16	: in std_logic := '0';
    B17	: in std_logic := '0';
    B18	: in std_logic := '0';

    C1	: in std_logic := '0';
    C2	: in std_logic := '0';
    C3	: in std_logic := '0';
    C4	: in std_logic := '0';
    C5	: in std_logic := '0';
    C6	: in std_logic := '0';
    C7	: in std_logic := '0';
    C8	: in std_logic := '0';
    C9	: in std_logic := '0';
    C10	: in std_logic := '0';
    C11	: in std_logic := '0';
    C12	: in std_logic := '0';
    C13	: in std_logic := '0';
    C14	: in std_logic := '0';
    C15	: in std_logic := '0';
    C16	: in std_logic := '0';
    C17	: in std_logic := '0';
    C18	: in std_logic := '0';
    C19	: in std_logic := '0';
    C20	: in std_logic := '0';
    C21	: in std_logic := '0';
    C22	: in std_logic := '0';
    C23	: in std_logic := '0';
    C24	: in std_logic := '0';
    C25	: in std_logic := '0';
    C26	: in std_logic := '0';
    C27	: in std_logic := '0';
    C28	: in std_logic := '0';
    C29	: in std_logic := '0';
    C30	: in std_logic := '0';
    C31	: in std_logic := '0';
    C32	: in std_logic := '0';
    C33	: in std_logic := '0';
    C34	: in std_logic := '0';
    C35	: in std_logic := '0';
    C36	: in std_logic := '0';

    CAI1	: in std_logic := '0';
    CAI2	: in std_logic := '0';
    CAI3	: in std_logic := '0';
    CAI4	: in std_logic := '0';
    CAI5	: in std_logic := '0';
    CAI6	: in std_logic := '0';
    CAI7	: in std_logic := '0';
    CAI8	: in std_logic := '0';
    CAI9	: in std_logic := '0';
    CAI10	: in std_logic := '0';
    CAI11	: in std_logic := '0';
    CAI12	: in std_logic := '0';
    CAI13	: in std_logic := '0';
    CAI14	: in std_logic := '0';
    CAI15	: in std_logic := '0';
    CAI16	: in std_logic := '0';
    CAI17	: in std_logic := '0';
    CAI18	: in std_logic := '0';
    CAI19	: in std_logic := '0';
    CAI20	: in std_logic := '0';
    CAI21	: in std_logic := '0';
    CAI22	: in std_logic := '0';
    CAI23	: in std_logic := '0';
    CAI24	: in std_logic := '0';

    CAO1	: out std_logic := '0';
    CAO2	: out std_logic := '0';
    CAO3	: out std_logic := '0';
    CAO4	: out std_logic := '0';
    CAO5	: out std_logic := '0';
    CAO6	: out std_logic := '0';
    CAO7	: out std_logic := '0';
    CAO8	: out std_logic := '0';
    CAO9	: out std_logic := '0';
    CAO10	: out std_logic := '0';
    CAO11	: out std_logic := '0';
    CAO12	: out std_logic := '0';
    CAO13	: out std_logic := '0';
    CAO14	: out std_logic := '0';
    CAO15	: out std_logic := '0';
    CAO16	: out std_logic := '0';
    CAO17	: out std_logic := '0';
    CAO18	: out std_logic := '0';
    CAO19	: out std_logic := '0';
    CAO20	: out std_logic := '0';
    CAO21	: out std_logic := '0';
    CAO22	: out std_logic := '0';
    CAO23	: out std_logic := '0';
    CAO24	: out std_logic := '0';

    CBI1	: in std_logic := '0';
    CBI2	: in std_logic := '0';
    CBI3	: in std_logic := '0';
    CBI4	: in std_logic := '0';
    CBI5	: in std_logic := '0';
    CBI6	: in std_logic := '0';
    CBI7	: in std_logic := '0';
    CBI8	: in std_logic := '0';
    CBI9	: in std_logic := '0';
    CBI10	: in std_logic := '0';
    CBI11	: in std_logic := '0';
    CBI12	: in std_logic := '0';
    CBI13	: in std_logic := '0';
    CBI14	: in std_logic := '0';
    CBI15	: in std_logic := '0';
    CBI16	: in std_logic := '0';
    CBI17	: in std_logic := '0';
    CBI18	: in std_logic := '0';

    CBO1	: out std_logic := '0';
    CBO2	: out std_logic := '0';
    CBO3	: out std_logic := '0';
    CBO4	: out std_logic := '0';
    CBO5	: out std_logic := '0';
    CBO6	: out std_logic := '0';
    CBO7	: out std_logic := '0';
    CBO8	: out std_logic := '0';
    CBO9	: out std_logic := '0';
    CBO10	: out std_logic := '0';
    CBO11	: out std_logic := '0';
    CBO12	: out std_logic := '0';
    CBO13	: out std_logic := '0';
    CBO14	: out std_logic := '0';
    CBO15	: out std_logic := '0';
    CBO16	: out std_logic := '0';
    CBO17	: out std_logic := '0';
    CBO18	: out std_logic := '0';

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO43	: out std_logic := '0';
    CO57	: out std_logic := '0';
    RESERVED	: out std_logic := '0';

    CZI1	: in std_logic := '0';
    CZI2	: in std_logic := '0';
    CZI3	: in std_logic := '0';
    CZI4	: in std_logic := '0';
    CZI5	: in std_logic := '0';
    CZI6	: in std_logic := '0';
    CZI7	: in std_logic := '0';
    CZI8	: in std_logic := '0';
    CZI9	: in std_logic := '0';
    CZI10	: in std_logic := '0';
    CZI11	: in std_logic := '0';
    CZI12	: in std_logic := '0';
    CZI13	: in std_logic := '0';
    CZI14	: in std_logic := '0';
    CZI15	: in std_logic := '0';
    CZI16	: in std_logic := '0';
    CZI17	: in std_logic := '0';
    CZI18	: in std_logic := '0';
    CZI19	: in std_logic := '0';
    CZI20	: in std_logic := '0';
    CZI21	: in std_logic := '0';
    CZI22	: in std_logic := '0';
    CZI23	: in std_logic := '0';
    CZI24	: in std_logic := '0';
    CZI25	: in std_logic := '0';
    CZI26	: in std_logic := '0';
    CZI27	: in std_logic := '0';
    CZI28	: in std_logic := '0';
    CZI29	: in std_logic := '0';
    CZI30	: in std_logic := '0';
    CZI31	: in std_logic := '0';
    CZI32	: in std_logic := '0';
    CZI33	: in std_logic := '0';
    CZI34	: in std_logic := '0';
    CZI35	: in std_logic := '0';
    CZI36	: in std_logic := '0';
    CZI37	: in std_logic := '0';
    CZI38	: in std_logic := '0';
    CZI39	: in std_logic := '0';
    CZI40	: in std_logic := '0';
    CZI41	: in std_logic := '0';
    CZI42	: in std_logic := '0';
    CZI43	: in std_logic := '0';
    CZI44	: in std_logic := '0';
    CZI45	: in std_logic := '0';
    CZI46	: in std_logic := '0';
    CZI47	: in std_logic := '0';
    CZI48	: in std_logic := '0';
    CZI49	: in std_logic := '0';
    CZI50	: in std_logic := '0';
    CZI51	: in std_logic := '0';
    CZI52	: in std_logic := '0';
    CZI53	: in std_logic := '0';
    CZI54	: in std_logic := '0';
    CZI55	: in std_logic := '0';
    CZI56	: in std_logic := '0';

    CZO1	: out std_logic := '0';
    CZO2	: out std_logic := '0';
    CZO3	: out std_logic := '0';
    CZO4	: out std_logic := '0';
    CZO5	: out std_logic := '0';
    CZO6	: out std_logic := '0';
    CZO7	: out std_logic := '0';
    CZO8	: out std_logic := '0';
    CZO9	: out std_logic := '0';
    CZO10	: out std_logic := '0';
    CZO11	: out std_logic := '0';
    CZO12	: out std_logic := '0';
    CZO13	: out std_logic := '0';
    CZO14	: out std_logic := '0';
    CZO15	: out std_logic := '0';
    CZO16	: out std_logic := '0';
    CZO17	: out std_logic := '0';
    CZO18	: out std_logic := '0';
    CZO19	: out std_logic := '0';
    CZO20	: out std_logic := '0';
    CZO21	: out std_logic := '0';
    CZO22	: out std_logic := '0';
    CZO23	: out std_logic := '0';
    CZO24	: out std_logic := '0';
    CZO25	: out std_logic := '0';
    CZO26	: out std_logic := '0';
    CZO27	: out std_logic := '0';
    CZO28	: out std_logic := '0';
    CZO29	: out std_logic := '0';
    CZO30	: out std_logic := '0';
    CZO31	: out std_logic := '0';
    CZO32	: out std_logic := '0';
    CZO33	: out std_logic := '0';
    CZO34	: out std_logic := '0';
    CZO35	: out std_logic := '0';
    CZO36	: out std_logic := '0';
    CZO37	: out std_logic := '0';
    CZO38	: out std_logic := '0';
    CZO39	: out std_logic := '0';
    CZO40	: out std_logic := '0';
    CZO41	: out std_logic := '0';
    CZO42	: out std_logic := '0';
    CZO43	: out std_logic := '0';
    CZO44	: out std_logic := '0';
    CZO45	: out std_logic := '0';
    CZO46	: out std_logic := '0';
    CZO47	: out std_logic := '0';
    CZO48	: out std_logic := '0';
    CZO49	: out std_logic := '0';
    CZO50	: out std_logic := '0';
    CZO51	: out std_logic := '0';
    CZO52	: out std_logic := '0';
    CZO53	: out std_logic := '0';
    CZO54	: out std_logic := '0';
    CZO55	: out std_logic := '0';
    CZO56	: out std_logic := '0';

    D1	: in std_logic := '0';
    D2	: in std_logic := '0';
    D3	: in std_logic := '0';
    D4	: in std_logic := '0';
    D5	: in std_logic := '0';
    D6	: in std_logic := '0';
    D7	: in std_logic := '0';
    D8	: in std_logic := '0';
    D9	: in std_logic := '0';
    D10	: in std_logic := '0';
    D11	: in std_logic := '0';
    D12	: in std_logic := '0';
    D13	: in std_logic := '0';
    D14	: in std_logic := '0';
    D15	: in std_logic := '0';
    D16	: in std_logic := '0';
    D17	: in std_logic := '0';
    D18	: in std_logic := '0';

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEZ	: in std_logic := '0';

    Z1	: out std_logic := '0';
    Z2	: out std_logic := '0';
    Z3	: out std_logic := '0';
    Z4	: out std_logic := '0';
    Z5	: out std_logic := '0';
    Z6	: out std_logic := '0';
    Z7	: out std_logic := '0';
    Z8	: out std_logic := '0';
    Z9	: out std_logic := '0';
    Z10	: out std_logic := '0';
    Z11	: out std_logic := '0';
    Z12	: out std_logic := '0';
    Z13	: out std_logic := '0';
    Z14	: out std_logic := '0';
    Z15	: out std_logic := '0';
    Z16	: out std_logic := '0';
    Z17	: out std_logic := '0';
    Z18	: out std_logic := '0';
    Z19	: out std_logic := '0';
    Z20	: out std_logic := '0';
    Z21	: out std_logic := '0';
    Z22	: out std_logic := '0';
    Z23	: out std_logic := '0';
    Z24	: out std_logic := '0';
    Z25	: out std_logic := '0';
    Z26	: out std_logic := '0';
    Z27	: out std_logic := '0';
    Z28	: out std_logic := '0';
    Z29	: out std_logic := '0';
    Z30	: out std_logic := '0';
    Z31	: out std_logic := '0';
    Z32	: out std_logic := '0';
    Z33	: out std_logic := '0';
    Z34	: out std_logic := '0';
    Z35	: out std_logic := '0';
    Z36	: out std_logic := '0';
    Z37	: out std_logic := '0';
    Z38	: out std_logic := '0';
    Z39	: out std_logic := '0';
    Z40	: out std_logic := '0';
    Z41	: out std_logic := '0';
    Z42	: out std_logic := '0';
    Z43	: out std_logic := '0';
    Z44	: out std_logic := '0';
    Z45	: out std_logic := '0';
    Z46	: out std_logic := '0';
    Z47	: out std_logic := '0';
    Z48	: out std_logic := '0';
    Z49	: out std_logic := '0';
    Z50	: out std_logic := '0';
    Z51	: out std_logic := '0';
    Z52	: out std_logic := '0';
    Z53	: out std_logic := '0';
    Z54	: out std_logic := '0';
    Z55	: out std_logic := '0';
    Z56	: out std_logic := '0'
    );
end component NX_DSP_U;

component NX_DSP_U_WRAP is
generic (
        std_mode    : string                  := "";
        raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
        raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
        raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
        raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
    );
port (
    A	: in std_logic_vector(23 downto 0) := (others => '0');
    B	: in std_logic_vector(17 downto 0) := (others => '0');
    C	: in std_logic_vector(35 downto 0) := (others => '0');

    CAI	: in std_logic_vector(23 downto 0) := (others => '0');
    CAO	: out std_logic_vector(23 downto 0) := (others => '0');
    CBI	: in std_logic_vector(17 downto 0) := (others => '0');
    CBO	: out std_logic_vector(17 downto 0) := (others => '0');

    CCI	: in std_logic := '0';
    CCO	: out std_logic := '0';
    CI	: in std_logic := '0';
    CK	: in std_logic := '0';
    CO43	: out std_logic := '0';
    CO57	: out std_logic := '0';

    CZI	: in std_logic_vector(55 downto 0) := (others => '0');
    CZO	: out std_logic_vector(55 downto 0) := (others => '0');

    D	: in std_logic_vector(17 downto 0) := (others => '0');

    OVF	: out std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEZ	: in std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0')
    );
end component NX_DSP_U_WRAP;

component NX_DSP_U_SPLIT is
generic (
        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
        ------------------------------------------------------------------------- 
        SIGNED_MODE        : bit                    := '0';
        INV_WE             : bit                    := '0';
        INV_WEZ            : bit                    := '0';
        INV_RST            : bit                    := '0';
        INV_RSTZ           : bit                    := '0';
        ALU_DYNAMIC_OP     : bit_vector(1 downto 0) := B"00";     -- "00" for Static,
        -- "-1" for Dynamic control from C
        -- "10" for Dynamic control from D
        SATURATION_RANK    : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB on Z and CZO result
        --(to define saturation and overflow)
        ENABLE_SATURATION  : bit                    := '0';       -- '0' for Disable,  '1' for Enable
        MUX_CCO            : bit                    := '0';       -- '0' for CC0 = ALU(42), '1' for CCO = ALU(56)
        MUX_Z              : bit                    := '0';       -- Select Z output. '0' for Y, '1' Saturation / ALU
        MUX_CZ             : bit                    := '0';       -- Select MUX_CZ input. '0' for CZI, '1' for CZO
        MUX_Y              : bit                    := '0';       -- Select ALU's Y input. '0' for MULT output, '1' for (B & A)
        MUX_X              : bit_vector(2 downto 0) := B"000";    -- Select MUX_X operation
        -- "000" for c[33:0]&d[41:34],
        -- "001" for C
        -- "010" for MUX_CZ[39:0]&C[15:0]
        -- "011" for MUX_CZ
        -- "100" for MUX_CZ >> 6
        -- "101" for MUX_CZ >> 12
        -- "110" for MUX_CZ >> 17
        -- "111" for MUX_CZ >> 18
        MUX_CCI            : bit                    := '0';       -- Select '1' input of CI mux. '0' for CCI, '1' for CO_feddback
        MUX_CI             : bit                    := '0';       -- Select input carry of ALU. '0' for CI, '1' for CCI/CO_feedback mux
        MUX_P              : bit                    := '0';       -- '1' for PRE_ADDER, '0' for B input
        MUX_B              : bit                    := '0';       -- '0' = B input, '1' = CBI input
        MUX_A              : bit                    := '0';       -- '0' = A input, '1' = CAI input
        PRE_ADDER_OP       : bit                    := '0';       -- '0' = Additon, '1' = Subraction

        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
        -------------------------------------------------------------------------
        PR_WE_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_WEZ_MUX         : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_RST_MUX         : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_RSTZ_MUX        : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_OV_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_CO_MUX          : bit                    := '0';       -- Registered carry out (CO42 & CO56)
        PR_CCO_MUX         : bit                    := '0';       -- Registered cascade carry out
        PR_Z_MUX           : bit                    := '0';       -- Registered output
        PR_CZ_MUX          : bit                    := '0';       -- Registered cascade output
        PR_Y_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_X_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_CI_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_MULT_MUX        : bit                    := '0';       -- No pipe reg  -- Register inside MULT
        PR_P_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
        PR_D_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_C_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_B_CASCADE_MUX   : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels for CAO output. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_B_MUX           : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels on B input. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_A_CASCADE_MUX   : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels for CAO output. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_A_MUX           : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels on A input. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
        -------------------------------------------------------------------------
        ENABLE_PR_OV_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CO_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CCO_RST  : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_Z_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CZ_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_Y_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_X_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CI_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_MULT_RST : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_P_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_D_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_C_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_B_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_A_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        -- PR_CZ_INIT         : bit_vector(5 downto 0) := B"000000"; -- Value of CZ's pipe register on reset

        -------------------------------------------------------------------------
        -- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
        -------------------------------------------------------------------------
        ALU_OP             : bit_vector(2 downto 0) := B"000"     -- ALU operation
        -- x+y+c    = "000"
        -- x-y-c    = "001"
        -- x-y+c-1  = "010"
        -- x+y-c+1  = "011"
        -- -x-y-c-1 = "100"
        -- -x+y+c-1 = "101"
        -- -x+y-c   = "110"
        -- -x-y+c-2 = "111"
    );
port (
    CK	: in std_logic := '0';
    R	: in std_logic := '0';
    RZ	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEZ	: in std_logic := '0';

    CI	: in std_logic := '0';
    A	: in std_logic_vector(23 downto 0) := (others => '0');
    B	: in std_logic_vector(17 downto 0) := (others => '0');
    C	: in std_logic_vector(35 downto 0) := (others => '0');
    D	: in std_logic_vector(17 downto 0) := (others => '0');
    CAI	: in std_logic_vector(23 downto 0) := (others => '0');
    CBI	: in std_logic_vector(17 downto 0) := (others => '0');
    CZI	: in std_logic_vector(55 downto 0) := (others => '0');
    CCI	: in std_logic := '0';

    Z	: out std_logic_vector(55 downto 0) := (others => '0');
    CO42	: out std_logic := '0';
    CO56	: out std_logic := '0';
    OVF	: out std_logic := '0';
    CAO	: out std_logic_vector(23 downto 0) := (others => '0');
    CBO	: out std_logic_vector(17 downto 0) := (others => '0');
    CZO	: out std_logic_vector(55 downto 0) := (others => '0');
    CCO	: out std_logic := '0'
    );
end component NX_DSP_U_SPLIT;

component NX_FIFO is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(5 downto 0) := "000000"
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    O	: out std_logic_vector(17 downto 0) := (others => '0');
    WRSTI	: in std_logic := '0';
    WAI	: in std_logic_vector(5 downto 0) := (others => '0');
    WAO	: out std_logic_vector(5 downto 0) := (others => '0');
    WEQ	: out std_logic := '0';
    RRSTI	: in std_logic := '0';
    RAI	: in std_logic_vector(5 downto 0) := (others => '0');
    RAO	: out std_logic_vector(5 downto 0) := (others => '0');
    REQ	: out std_logic := '0'
);
end component NX_FIFO;

component NX_XFIFO_64x18 is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    O	: out std_logic_vector(17 downto 0) := (others => '0');
    WRSTI	: in std_logic := '0';
    WAI	: in std_logic_vector(6 downto 0) := (others => '0');
    WAO	: out std_logic_vector(6 downto 0) := (others => '0');
    WEQ	: out std_logic_vector(1 downto 0) := (others => '0');
    RRSTI	: in std_logic := '0';
    RAI	: in std_logic_vector(6 downto 0) := (others => '0');
    RAO	: out std_logic_vector(6 downto 0) := (others => '0');
    REQ	: out std_logic_vector(1 downto 0) := (others => '0')
);
end component NX_XFIFO_64x18;

component NX_XFIFO_32x36 is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0';
    I	: in std_logic_vector(35 downto 0) := (others => '0');
    O	: out std_logic_vector(35 downto 0) := (others => '0');
    WRSTI	: in std_logic := '0';
    WAI	: in std_logic_vector(5 downto 0) := (others => '0');
    WAO	: out std_logic_vector(5 downto 0) := (others => '0');
    WEQ	: out std_logic := '0';
    RRSTI	: in std_logic := '0';
    RAI	: in std_logic_vector(5 downto 0) := (others => '0');
    RAO	: out std_logic_vector(5 downto 0) := (others => '0');
    REQ	: out std_logic := '0'
);
end component NX_XFIFO_32x36;

component NX_FIFO_U is
generic (
    mode           : integer := 0; -- 0: DPREG - 1: XFIFO_64x18 - 2: XFIFO_32x36
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0';
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    I5	: in std_logic := '0';
    I6	: in std_logic := '0';
    I7	: in std_logic := '0';
    I8	: in std_logic := '0';
    I9	: in std_logic := '0';
    I10	: in std_logic := '0';
    I11	: in std_logic := '0';
    I12	: in std_logic := '0';
    I13	: in std_logic := '0';
    I14	: in std_logic := '0';
    I15	: in std_logic := '0';
    I16	: in std_logic := '0';
    I17	: in std_logic := '0';
    I18	: in std_logic := '0';
    I19	: in std_logic := '0';
    I20	: in std_logic := '0';
    I21	: in std_logic := '0';
    I22	: in std_logic := '0';
    I23	: in std_logic := '0';
    I24	: in std_logic := '0';
    I25	: in std_logic := '0';
    I26	: in std_logic := '0';
    I27	: in std_logic := '0';
    I28	: in std_logic := '0';
    I29	: in std_logic := '0';
    I30	: in std_logic := '0';
    I31	: in std_logic := '0';
    I32	: in std_logic := '0';
    I33	: in std_logic := '0';
    I34	: in std_logic := '0';
    I35	: in std_logic := '0';
    I36	: in std_logic := '0';
    O1	: out std_logic := '0';
    O2	: out std_logic := '0';
    O3	: out std_logic := '0';
    O4	: out std_logic := '0';
    O5	: out std_logic := '0';
    O6	: out std_logic := '0';
    O7	: out std_logic := '0';
    O8	: out std_logic := '0';
    O9	: out std_logic := '0';
    O10	: out std_logic := '0';
    O11	: out std_logic := '0';
    O12	: out std_logic := '0';
    O13	: out std_logic := '0';
    O14	: out std_logic := '0';
    O15	: out std_logic := '0';
    O16	: out std_logic := '0';
    O17	: out std_logic := '0';
    O18	: out std_logic := '0';
    O19	: out std_logic := '0';
    O20	: out std_logic := '0';
    O21	: out std_logic := '0';
    O22	: out std_logic := '0';
    O23	: out std_logic := '0';
    O24	: out std_logic := '0';
    O25	: out std_logic := '0';
    O26	: out std_logic := '0';
    O27	: out std_logic := '0';
    O28	: out std_logic := '0';
    O29	: out std_logic := '0';
    O30	: out std_logic := '0';
    O31	: out std_logic := '0';
    O32	: out std_logic := '0';
    O33	: out std_logic := '0';
    O34	: out std_logic := '0';
    O35	: out std_logic := '0';
    O36	: out std_logic := '0';
    WRSTI	: in std_logic := '0';
    WAI1	: in std_logic := '0';
    WAI2	: in std_logic := '0';
    WAI3	: in std_logic := '0';
    WAI4	: in std_logic := '0';
    WAI5	: in std_logic := '0';
    WAI6	: in std_logic := '0';
    WAI7	: in std_logic := '0';
    WAO1	: out std_logic := '0';
    WAO2	: out std_logic := '0';
    WAO3	: out std_logic := '0';
    WAO4	: out std_logic := '0';
    WAO5	: out std_logic := '0';
    WAO6	: out std_logic := '0';
    WAO7	: out std_logic := '0';
    WEQ1	: out std_logic := '0';
    WEQ2	: out std_logic := '0';
    RRSTI	: in std_logic := '0';
    RAI1	: in std_logic := '0';
    RAI2	: in std_logic := '0';
    RAI3	: in std_logic := '0';
    RAI4	: in std_logic := '0';
    RAI5	: in std_logic := '0';
    RAI6	: in std_logic := '0';
    RAI7	: in std_logic := '0';
    RAO1	: out std_logic := '0';
    RAO2	: out std_logic := '0';
    RAO3	: out std_logic := '0';
    RAO4	: out std_logic := '0';
    RAO5	: out std_logic := '0';
    RAO6	: out std_logic := '0';
    RAO7	: out std_logic := '0';
    REQ1	: out std_logic := '0';
    REQ2	: out std_logic := '0'
);
end component NX_FIFO_U;

component NX_GCK_U is
generic (
    inv_in   : bit    := '0';
    inv_out  : bit    := '0';
    std_mode : string := "BYPASS" -- MUX / CKS / BYPASS / CSC
);
port (
    SI1	: in std_logic := '0';
    SI2	: in std_logic := '0';
    CMD	: in std_logic := '0';
    SO	: out std_logic := '0'
);
end component NX_GCK_U;

component NX_CRX_L is
generic (
     test                         : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc           : bit := '0';
     pcs_bypass_usr_cdc           : bit := '0';
     pcs_debug_en                 : bit := '0';
     pcs_fsm_watchdog_en          : bit := '0';
     pma_clk_pos                  : bit := '0';
     pcs_protocol_size            : bit := '0';
     pcs_loopback                 : bit := '0';
     pcs_polarity                 : bit := '0';
     pcs_p_comma_en               : bit := '0';
     pcs_p_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_m_comma_en               : bit := '0';
     pcs_m_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_comma_mask               : bit_vector(9 downto 0) := (others => '0');
     pcs_nb_comma_bef_realign     : bit_vector(1 downto 0) := (others => '0');
     pcs_align_bypass             : bit := '0';
     pcs_dec_bypass               : bit := '0';
     pcs_el_buff_max_comp         : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_diff_bef_comp    : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_only_one_skp     : bit := '0';
     pcs_el_buff_underflow_handle : bit := '0';
     pcs_el_buff_skp_seq_size     : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_char_0       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_1       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_2       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_3       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_size  : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_header_0     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_1     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_2     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_3     : bit_vector(8 downto 0) := (others => '0');
     pcs_buffers_use_cdc          : bit := '0';
     pcs_buffers_bypass           : bit := '0';
     pcs_sync_supported           : bit := '0';
     pcs_replace_bypass           : bit := '0';
     pcs_dscr_bypass              : bit := '0';
     pcs_8b_dscr_sel              : bit := '0';
     pcs_fsm_sel                  : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divf_en_n            : bit := '0';
     pma_pll_divm_en_n            : bit := '0';
     pma_pll_divn_en_n            : bit := '0';
     pma_cdr_cp                   : bit_vector(3 downto 0) := (others => '0');
     pma_ctrl_term                : bit_vector(5 downto 0) := (others => '0');
     pma_pll_cpump_n              : bit_vector(2 downto 0) := (others => '0');
     pma_pll_divf                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divm                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divn                 : bit := '0';
     pma_loopback                 : bit := '0';
     location                     : string := ""
 );
port (
    DSCR_E_I	: in std_logic := '0';
    DEC_E_I	: in std_logic := '0';
    ALIGN_E_I	: in std_logic := '0';
    ALIGN_S_I	: in std_logic := '0';
    REP_E_I	: in std_logic := '0';
    BUF_R_I	: in std_logic := '0';

    OVS_BS_I1	: in std_logic := '0';
    OVS_BS_I2	: in std_logic := '0';

    BUF_FE_I	: in std_logic := '0';
    RST_N_I	: in std_logic := '0';
    CDR_R_I	: in std_logic := '0';
    CKG_RN_I	: in std_logic := '0';
    PLL_RN_I	: in std_logic := '0';

    TST_I1	: in std_logic := '0';
    TST_I2	: in std_logic := '0';
    TST_I3	: in std_logic := '0';
    TST_I4	: in std_logic := '0';

    LOS_O	: out std_logic := '0';

    DATA_O1	: out std_logic := '0';
    DATA_O2	: out std_logic := '0';
    DATA_O3	: out std_logic := '0';
    DATA_O4	: out std_logic := '0';
    DATA_O5	: out std_logic := '0';
    DATA_O6	: out std_logic := '0';
    DATA_O7	: out std_logic := '0';
    DATA_O8	: out std_logic := '0';
    DATA_O9	: out std_logic := '0';
    DATA_O10	: out std_logic := '0';
    DATA_O11	: out std_logic := '0';
    DATA_O12	: out std_logic := '0';
    DATA_O13	: out std_logic := '0';
    DATA_O14	: out std_logic := '0';
    DATA_O15	: out std_logic := '0';
    DATA_O16	: out std_logic := '0';
    DATA_O17	: out std_logic := '0';
    DATA_O18	: out std_logic := '0';
    DATA_O19	: out std_logic := '0';
    DATA_O20	: out std_logic := '0';
    DATA_O21	: out std_logic := '0';
    DATA_O22	: out std_logic := '0';
    DATA_O23	: out std_logic := '0';
    DATA_O24	: out std_logic := '0';
    DATA_O25	: out std_logic := '0';
    DATA_O26	: out std_logic := '0';
    DATA_O27	: out std_logic := '0';
    DATA_O28	: out std_logic := '0';
    DATA_O29	: out std_logic := '0';
    DATA_O30	: out std_logic := '0';
    DATA_O31	: out std_logic := '0';
    DATA_O32	: out std_logic := '0';
    DATA_O33	: out std_logic := '0';
    DATA_O34	: out std_logic := '0';
    DATA_O35	: out std_logic := '0';
    DATA_O36	: out std_logic := '0';
    DATA_O37	: out std_logic := '0';
    DATA_O38	: out std_logic := '0';
    DATA_O39	: out std_logic := '0';
    DATA_O40	: out std_logic := '0';
    DATA_O41	: out std_logic := '0';
    DATA_O42	: out std_logic := '0';
    DATA_O43	: out std_logic := '0';
    DATA_O44	: out std_logic := '0';
    DATA_O45	: out std_logic := '0';
    DATA_O46	: out std_logic := '0';
    DATA_O47	: out std_logic := '0';
    DATA_O48	: out std_logic := '0';
    DATA_O49	: out std_logic := '0';
    DATA_O50	: out std_logic := '0';
    DATA_O51	: out std_logic := '0';
    DATA_O52	: out std_logic := '0';
    DATA_O53	: out std_logic := '0';
    DATA_O54	: out std_logic := '0';
    DATA_O55	: out std_logic := '0';
    DATA_O56	: out std_logic := '0';
    DATA_O57	: out std_logic := '0';
    DATA_O58	: out std_logic := '0';
    DATA_O59	: out std_logic := '0';
    DATA_O60	: out std_logic := '0';
    DATA_O61	: out std_logic := '0';
    DATA_O62	: out std_logic := '0';
    DATA_O63	: out std_logic := '0';
    DATA_O64	: out std_logic := '0';

    CH_COM_O1	: out std_logic := '0';
    CH_COM_O2	: out std_logic := '0';
    CH_COM_O3	: out std_logic := '0';
    CH_COM_O4	: out std_logic := '0';
    CH_COM_O5	: out std_logic := '0';
    CH_COM_O6	: out std_logic := '0';
    CH_COM_O7	: out std_logic := '0';
    CH_COM_O8	: out std_logic := '0';

    CH_K_O1	: out std_logic := '0';
    CH_K_O2	: out std_logic := '0';
    CH_K_O3	: out std_logic := '0';
    CH_K_O4	: out std_logic := '0';
    CH_K_O5	: out std_logic := '0';
    CH_K_O6	: out std_logic := '0';
    CH_K_O7	: out std_logic := '0';
    CH_K_O8	: out std_logic := '0';

    NIT_O1	: out std_logic := '0';
    NIT_O2	: out std_logic := '0';
    NIT_O3	: out std_logic := '0';
    NIT_O4	: out std_logic := '0';
    NIT_O5	: out std_logic := '0';
    NIT_O6	: out std_logic := '0';
    NIT_O7	: out std_logic := '0';
    NIT_O8	: out std_logic := '0';

    D_ERR_O1	: out std_logic := '0';
    D_ERR_O2	: out std_logic := '0';
    D_ERR_O3	: out std_logic := '0';
    D_ERR_O4	: out std_logic := '0';
    D_ERR_O5	: out std_logic := '0';
    D_ERR_O6	: out std_logic := '0';
    D_ERR_O7	: out std_logic := '0';
    D_ERR_O8	: out std_logic := '0';

    CH_A_O1	: out std_logic := '0';
    CH_A_O2	: out std_logic := '0';
    CH_A_O3	: out std_logic := '0';
    CH_A_O4	: out std_logic := '0';
    CH_A_O5	: out std_logic := '0';
    CH_A_O6	: out std_logic := '0';
    CH_A_O7	: out std_logic := '0';
    CH_A_O8	: out std_logic := '0';

    CH_F_O1	: out std_logic := '0';
    CH_F_O2	: out std_logic := '0';
    CH_F_O3	: out std_logic := '0';
    CH_F_O4	: out std_logic := '0';
    CH_F_O5	: out std_logic := '0';
    CH_F_O6	: out std_logic := '0';
    CH_F_O7	: out std_logic := '0';
    CH_F_O8	: out std_logic := '0';

    ALIGN_O	: out std_logic := '0';
    BUSY_O	: out std_logic := '0';

    TST_O1	: out std_logic := '0';
    TST_O2	: out std_logic := '0';
    TST_O3	: out std_logic := '0';
    TST_O4	: out std_logic := '0';
    TST_O5	: out std_logic := '0';
    TST_O6	: out std_logic := '0';
    TST_O7	: out std_logic := '0';
    TST_O8	: out std_logic := '0';

    LOCK_O	: out std_logic := '0';

    LINK	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');

    RX_I	: in std_logic := '0'
);
end component NX_CRX_L;

component NX_CTX_L is
generic (
     pma_clk_pos          : bit := '0';
     pcs_protocol_size    : bit := '0';
     pcs_8b_scr_sel       : bit := '0';
     pcs_scr_init         : bit_vector(16 downto 0) := (others => '0');
     pcs_scr_bypass       : bit := '0';
     pcs_sync_supported   : bit := '0';
     pcs_replace_bypass   : bit := '0';
     pcs_enc_bypass       : bit := '0';
     pcs_loopback         : bit := '0';
     pcs_polarity         : bit := '0';
     pcs_esistream_fsm_en : bit := '0';
     test                 : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc   : bit := '0';
     pcs_bypass_usr_cdc   : bit := '0';
     pma_loopback         : bit := '0';
     location             : string := ""
 );
port (
    ENC_E_I1	: in std_logic := '0';
    ENC_E_I2	: in std_logic := '0';
    ENC_E_I3	: in std_logic := '0';
    ENC_E_I4	: in std_logic := '0';
    ENC_E_I5	: in std_logic := '0';
    ENC_E_I6	: in std_logic := '0';
    ENC_E_I7	: in std_logic := '0';
    ENC_E_I8	: in std_logic := '0';

    CH_K_I1	: in std_logic := '0';
    CH_K_I2	: in std_logic := '0';
    CH_K_I3	: in std_logic := '0';
    CH_K_I4	: in std_logic := '0';
    CH_K_I5	: in std_logic := '0';
    CH_K_I6	: in std_logic := '0';
    CH_K_I7	: in std_logic := '0';
    CH_K_I8	: in std_logic := '0';

    SCR_E_I1	: in std_logic := '0';
    SCR_E_I2	: in std_logic := '0';
    SCR_E_I3	: in std_logic := '0';
    SCR_E_I4	: in std_logic := '0';
    SCR_E_I5	: in std_logic := '0';
    SCR_E_I6	: in std_logic := '0';
    SCR_E_I7	: in std_logic := '0';
    SCR_E_I8	: in std_logic := '0';

    EOMF_I1	: in std_logic := '0';
    EOMF_I2	: in std_logic := '0';
    EOMF_I3	: in std_logic := '0';
    EOMF_I4	: in std_logic := '0';
    EOMF_I5	: in std_logic := '0';
    EOMF_I6	: in std_logic := '0';
    EOMF_I7	: in std_logic := '0';
    EOMF_I8	: in std_logic := '0';

    EOF_I1	: in std_logic := '0';
    EOF_I2	: in std_logic := '0';
    EOF_I3	: in std_logic := '0';
    EOF_I4	: in std_logic := '0';
    EOF_I5	: in std_logic := '0';
    EOF_I6	: in std_logic := '0';
    EOF_I7	: in std_logic := '0';
    EOF_I8	: in std_logic := '0';

    REP_E_I	: in std_logic := '0';
    RST_N_I	: in std_logic := '0';

    TST_I1	: in std_logic := '0';
    TST_I2	: in std_logic := '0';
    TST_I3	: in std_logic := '0';
    TST_I4	: in std_logic := '0';

    DATA_I1	: in std_logic := '0';
    DATA_I2	: in std_logic := '0';
    DATA_I3	: in std_logic := '0';
    DATA_I4	: in std_logic := '0';
    DATA_I5	: in std_logic := '0';
    DATA_I6	: in std_logic := '0';
    DATA_I7	: in std_logic := '0';
    DATA_I8	: in std_logic := '0';
    DATA_I9	: in std_logic := '0';
    DATA_I10	: in std_logic := '0';
    DATA_I11	: in std_logic := '0';
    DATA_I12	: in std_logic := '0';
    DATA_I13	: in std_logic := '0';
    DATA_I14	: in std_logic := '0';
    DATA_I15	: in std_logic := '0';
    DATA_I16	: in std_logic := '0';
    DATA_I17	: in std_logic := '0';
    DATA_I18	: in std_logic := '0';
    DATA_I19	: in std_logic := '0';
    DATA_I20	: in std_logic := '0';
    DATA_I21	: in std_logic := '0';
    DATA_I22	: in std_logic := '0';
    DATA_I23	: in std_logic := '0';
    DATA_I24	: in std_logic := '0';
    DATA_I25	: in std_logic := '0';
    DATA_I26	: in std_logic := '0';
    DATA_I27	: in std_logic := '0';
    DATA_I28	: in std_logic := '0';
    DATA_I29	: in std_logic := '0';
    DATA_I30	: in std_logic := '0';
    DATA_I31	: in std_logic := '0';
    DATA_I32	: in std_logic := '0';
    DATA_I33	: in std_logic := '0';
    DATA_I34	: in std_logic := '0';
    DATA_I35	: in std_logic := '0';
    DATA_I36	: in std_logic := '0';
    DATA_I37	: in std_logic := '0';
    DATA_I38	: in std_logic := '0';
    DATA_I39	: in std_logic := '0';
    DATA_I40	: in std_logic := '0';
    DATA_I41	: in std_logic := '0';
    DATA_I42	: in std_logic := '0';
    DATA_I43	: in std_logic := '0';
    DATA_I44	: in std_logic := '0';
    DATA_I45	: in std_logic := '0';
    DATA_I46	: in std_logic := '0';
    DATA_I47	: in std_logic := '0';
    DATA_I48	: in std_logic := '0';
    DATA_I49	: in std_logic := '0';
    DATA_I50	: in std_logic := '0';
    DATA_I51	: in std_logic := '0';
    DATA_I52	: in std_logic := '0';
    DATA_I53	: in std_logic := '0';
    DATA_I54	: in std_logic := '0';
    DATA_I55	: in std_logic := '0';
    DATA_I56	: in std_logic := '0';
    DATA_I57	: in std_logic := '0';
    DATA_I58	: in std_logic := '0';
    DATA_I59	: in std_logic := '0';
    DATA_I60	: in std_logic := '0';
    DATA_I61	: in std_logic := '0';
    DATA_I62	: in std_logic := '0';
    DATA_I63	: in std_logic := '0';
    DATA_I64	: in std_logic := '0';

    TST_O1	: out std_logic := '0';
    TST_O2	: out std_logic := '0';
    TST_O3	: out std_logic := '0';
    TST_O4	: out std_logic := '0';

    BUSY_O	: out std_logic := '0';
    CLK_E_I	: in std_logic := '0';

    LINK	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');

    TX_O	: out std_logic := '0'
);
end component NX_CTX_L;

component NX_HSSL_L_FULL is
generic (
   cfg_main_i : bit_vector( 33 downto 0) := (others => '0');
   cfg_tx0_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx0_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx1_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx1_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx2_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx2_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx3_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx3_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx4_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx4_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx5_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx5_i  : bit_vector(159 downto 0) := (others => '0');
   location   : string := ""
 );
port (
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ MAIN ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- Fabric Interface
    hssl_clk_user_i	: in std_logic := '0';
    hssl_clk_ref_i	: in std_logic := '0';
    hssl_clock_o	: out std_logic := '0';
    usr_com_tx_pma_pre_sign_i	: in std_logic := '0';
    usr_com_tx_pma_pre_en_i	: in std_logic := '0';
    usr_com_tx_pma_pre_input_sel_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_tx_pma_main_sign_i	: in std_logic := '0';
    usr_com_rx_pma_m_eye_i	: in std_logic := '0';
    usr_com_tx_pma_main_en_i	: in std_logic_vector(5 downto 0) := (others => '0');
    usr_com_tx_pma_margin_sel_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_tx_pma_margin_input_sel_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_tx_pma_margin_sel_var_i	: in std_logic_vector(4 downto 0) := (others => '0');
    usr_com_tx_pma_margin_input_sel_var_i	: in std_logic_vector(4 downto 0) := (others => '0');
    usr_com_tx_pma_post_en_i	: in std_logic_vector(4 downto 0) := (others => '0');
    usr_com_tx_pma_post_sign_i	: in std_logic := '0';
    usr_com_tx_pma_post_input_sel_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_tx_pma_post_input_sel_var_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_rx_pma_ctle_cap_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_rx_pma_ctle_resp_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_rx_pma_ctle_resn_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_com_ctrl_tx_sel_i	: in std_logic_vector(5 downto 0) := (others => '0');
    usr_com_ctrl_rx_sel_i	: in std_logic_vector(5 downto 0) := (others => '0');
    usr_pll_pma_rst_n_i	: in std_logic := '0';
    usr_main_rst_n_i	: in std_logic := '0';
    usr_calibrate_pma_res_p1_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_calibrate_pma_res_n2_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_calibrate_pma_res_n3_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_calibrate_pma_res_p4_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_calibrate_pma_sel_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_calibrate_pma_en_i	: in std_logic := '0';
    usr_pcs_ctrl_pll_lock_en_i	: in std_logic := '0';
    usr_pcs_ctrl_ovs_en_i	: in std_logic := '0';
    usr_main_test_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_pll_lock_o	: out std_logic := '0';
    usr_calibrate_pma_out_o	: out std_logic := '0';
    usr_main_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    pma_clk_ext_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 0 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx0_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx0_rst_n_i	: in std_logic := '0';
    usr_tx0_pma_clk_en_i	: in std_logic := '0';
    usr_tx0_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx0_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx0_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx0_busy_o	: out std_logic := '0';
    pma_tx0_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx0_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx0_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx0_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx0_ctrl_align_en_i	: in std_logic := '0';
    usr_rx0_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx0_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx0_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx0_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx0_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx0_rst_n_i	: in std_logic := '0';
    usr_rx0_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx0_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx0_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx0_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx0_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx0_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx0_busy_o	: out std_logic := '0';
    usr_rx0_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_pll_lock_o	: out std_logic := '0';
    pma_rx0_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 1 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx1_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx1_rst_n_i	: in std_logic := '0';
    usr_tx1_pma_clk_en_i	: in std_logic := '0';
    usr_tx1_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx1_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx1_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx1_busy_o	: out std_logic := '0';
    pma_tx1_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx1_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx1_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx1_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx1_ctrl_align_en_i	: in std_logic := '0';
    usr_rx1_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx1_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx1_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx1_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx1_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx1_rst_n_i	: in std_logic := '0';
    usr_rx1_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx1_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx1_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx1_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx1_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx1_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx1_busy_o	: out std_logic := '0';
    usr_rx1_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_pll_lock_o	: out std_logic := '0';
    pma_rx1_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 2 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx2_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx2_rst_n_i	: in std_logic := '0';
    usr_tx2_pma_clk_en_i	: in std_logic := '0';
    usr_tx2_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx2_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx2_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx2_busy_o	: out std_logic := '0';
    pma_tx2_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx2_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx2_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx2_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx2_ctrl_align_en_i	: in std_logic := '0';
    usr_rx2_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx2_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx2_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx2_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx2_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx2_rst_n_i	: in std_logic := '0';
    usr_rx2_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx2_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx2_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx2_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx2_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx2_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx2_busy_o	: out std_logic := '0';
    usr_rx2_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_pll_lock_o	: out std_logic := '0';
    pma_rx2_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 3 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx3_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx3_rst_n_i	: in std_logic := '0';
    usr_tx3_pma_clk_en_i	: in std_logic := '0';
    usr_tx3_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx3_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx3_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx3_busy_o	: out std_logic := '0';
    pma_tx3_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx3_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx3_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx3_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx3_ctrl_align_en_i	: in std_logic := '0';
    usr_rx3_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx3_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx3_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx3_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx3_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx3_rst_n_i	: in std_logic := '0';
    usr_rx3_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx3_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx3_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx3_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx3_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx3_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx3_busy_o	: out std_logic := '0';
    usr_rx3_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_pll_lock_o	: out std_logic := '0';
    pma_rx3_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 4 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx4_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx4_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx4_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx4_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx4_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx4_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx4_rst_n_i	: in std_logic := '0';
    usr_tx4_pma_clk_en_i	: in std_logic := '0';
    usr_tx4_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx4_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx4_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx4_busy_o	: out std_logic := '0';
    pma_tx4_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx4_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx4_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx4_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx4_ctrl_align_en_i	: in std_logic := '0';
    usr_rx4_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx4_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx4_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx4_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx4_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx4_rst_n_i	: in std_logic := '0';
    usr_rx4_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx4_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx4_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx4_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx4_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx4_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx4_busy_o	: out std_logic := '0';
    usr_rx4_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx4_pll_lock_o	: out std_logic := '0';
    pma_rx4_i	: in std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 5 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
    usr_tx5_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx5_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx5_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx5_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx5_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx5_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx5_rst_n_i	: in std_logic := '0';
    usr_tx5_pma_clk_en_i	: in std_logic := '0';
    usr_tx5_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_tx5_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx5_test_o	: out std_logic_vector(3 downto 0) := (others => '0');
    usr_tx5_busy_o	: out std_logic := '0';
    pma_tx5_o	: out std_logic := '0';
    -- RX - Fabric Interface
    usr_rx5_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx5_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx5_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx5_ctrl_align_en_i	: in std_logic := '0';
    usr_rx5_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx5_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx5_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx5_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx5_ctrl_el_buff_fifo_en_i	: in std_logic := '0';
    usr_rx5_rst_n_i	: in std_logic := '0';
    usr_rx5_pma_cdr_rst_i	: in std_logic := '0';
    usr_rx5_pma_ckgen_rst_n_i	: in std_logic := '0';
    usr_rx5_pma_pll_rst_n_i	: in std_logic := '0';
    usr_rx5_test_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_rx5_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx5_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx5_busy_o	: out std_logic := '0';
    usr_rx5_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx5_pll_lock_o	: out std_logic := '0';
    pma_rx5_i	: in std_logic := '0'
);
end component NX_HSSL_L_FULL;

component NX_PMA_L is
generic (
     main_test                   : bit_vector(7 downto 0) := (others => '0');
     rx_pma_half_step            : bit := '0';
     pll_pma_int_data_len        : bit := '0';
     pll_pma_cpump_n             : bit_vector(2 downto 0) := (others => '0');
     pll_pma_divf                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divm                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divn                : bit := '0';
     pll_pma_lvds_mux            : bit := '0';
     pll_pma_mux_ckref           : bit := '0';
     pll_pma_divf_en_n           : bit := '0';
     pll_pma_divm_en_n           : bit := '0';
     pll_pma_divn_en_n           : bit := '0';
     main_clk_to_fabric_div_mode : bit := '0';
     main_clk_to_fabric_div_en   : bit := '0';
     main_clk_to_fabric_sel      : bit := '0';
     main_use_only_usr_clock     : bit := '0';
     main_use_pcs_clk_2          : bit := '0';
     pcs_word_len                : bit_vector(1 downto 0) := (others => '0');
     pcs_ovs_mode                : bit := '0';
     pcs_pll_lock_count          : bit_vector(2 downto 0) := (others => '0');
     location                    : string := ""
 );
port (
    CLK_USER_I	: in std_logic := '0';
    CLK_REF_I	: in std_logic := '0';
--    CLK_I1      : in  std_logic;
--    CLK_I2      : in  std_logic;
--    CLK_I3      : in  std_logic;
--    CLK_I4      : in  std_logic;
--    CLK_I5      : in  std_logic;
--    CLK_I6      : in  std_logic;
--    CLK_I7      : in  std_logic;
--    CLK_I8      : in  std_logic;

    PRE_SG_I	: in std_logic := '0';
    PRE_EN_I	: in std_logic := '0';

    PRE_IS_I1	: in std_logic := '0';
    PRE_IS_I2	: in std_logic := '0';
    PRE_IS_I3	: in std_logic := '0';
    PRE_IS_I4	: in std_logic := '0';

    MAIN_SG_I	: in std_logic := '0';

    MAIN_EN_I1	: in std_logic := '0';
    MAIN_EN_I2	: in std_logic := '0';
    MAIN_EN_I3	: in std_logic := '0';
    MAIN_EN_I4	: in std_logic := '0';
    MAIN_EN_I5	: in std_logic := '0';
    MAIN_EN_I6	: in std_logic := '0';

    MARG_S_I1	: in std_logic := '0';
    MARG_S_I2	: in std_logic := '0';
    MARG_S_I3	: in std_logic := '0';
    MARG_S_I4	: in std_logic := '0';

    MARG_IS_I1	: in std_logic := '0';
    MARG_IS_I2	: in std_logic := '0';
    MARG_IS_I3	: in std_logic := '0';
    MARG_IS_I4	: in std_logic := '0';

    MARG_SV_I1	: in std_logic := '0';
    MARG_SV_I2	: in std_logic := '0';
    MARG_SV_I3	: in std_logic := '0';
    MARG_SV_I4	: in std_logic := '0';
    MARG_SV_I5	: in std_logic := '0';

    MARG_ISV_I1	: in std_logic := '0';
    MARG_ISV_I2	: in std_logic := '0';
    MARG_ISV_I3	: in std_logic := '0';
    MARG_ISV_I4	: in std_logic := '0';
    MARG_ISV_I5	: in std_logic := '0';

    POST_EN_I1	: in std_logic := '0';
    POST_EN_I2	: in std_logic := '0';
    POST_EN_I3	: in std_logic := '0';
    POST_EN_I4	: in std_logic := '0';
    POST_EN_I5	: in std_logic := '0';

    POST_SG_I	: in std_logic := '0';

    POST_IS_I1	: in std_logic := '0';
    POST_IS_I2	: in std_logic := '0';
    POST_IS_I3	: in std_logic := '0';
    POST_IS_I4	: in std_logic := '0';

    POST_ISV_I1	: in std_logic := '0';
    POST_ISV_I2	: in std_logic := '0';
    POST_ISV_I3	: in std_logic := '0';
    POST_ISV_I4	: in std_logic := '0';

    TX_SEL_I1	: in std_logic := '0';
    TX_SEL_I2	: in std_logic := '0';
    TX_SEL_I3	: in std_logic := '0';
    TX_SEL_I4	: in std_logic := '0';
    TX_SEL_I5	: in std_logic := '0';
    TX_SEL_I6	: in std_logic := '0';

    CT_CAP_I1	: in std_logic := '0';
    CT_CAP_I2	: in std_logic := '0';
    CT_CAP_I3	: in std_logic := '0';
    CT_CAP_I4	: in std_logic := '0';

    CT_RESP_I1	: in std_logic := '0';
    CT_RESP_I2	: in std_logic := '0';
    CT_RESP_I3	: in std_logic := '0';
    CT_RESP_I4	: in std_logic := '0';

    CT_RESN_I1	: in std_logic := '0';
    CT_RESN_I2	: in std_logic := '0';
    CT_RESN_I3	: in std_logic := '0';
    CT_RESN_I4	: in std_logic := '0';

    M_EYE_I	: in std_logic := '0';

    RX_SEL_I1	: in std_logic := '0';
    RX_SEL_I2	: in std_logic := '0';
    RX_SEL_I3	: in std_logic := '0';
    RX_SEL_I4	: in std_logic := '0';
    RX_SEL_I5	: in std_logic := '0';
    RX_SEL_I6	: in std_logic := '0';

    PLL_RN_I	: in std_logic := '0';
    RST_N_I	: in std_logic := '0';

    CAL_1P_I1	: in std_logic := '0';
    CAL_1P_I2	: in std_logic := '0';
    CAL_1P_I3	: in std_logic := '0';
    CAL_1P_I4	: in std_logic := '0';
    CAL_1P_I5	: in std_logic := '0';
    CAL_1P_I6	: in std_logic := '0';
    CAL_1P_I7	: in std_logic := '0';
    CAL_1P_I8	: in std_logic := '0';

    CAL_2N_I1	: in std_logic := '0';
    CAL_2N_I2	: in std_logic := '0';
    CAL_2N_I3	: in std_logic := '0';
    CAL_2N_I4	: in std_logic := '0';
    CAL_2N_I5	: in std_logic := '0';
    CAL_2N_I6	: in std_logic := '0';
    CAL_2N_I7	: in std_logic := '0';
    CAL_2N_I8	: in std_logic := '0';

    CAL_3N_I1	: in std_logic := '0';
    CAL_3N_I2	: in std_logic := '0';
    CAL_3N_I3	: in std_logic := '0';
    CAL_3N_I4	: in std_logic := '0';
    CAL_3N_I5	: in std_logic := '0';
    CAL_3N_I6	: in std_logic := '0';
    CAL_3N_I7	: in std_logic := '0';
    CAL_3N_I8	: in std_logic := '0';

    CAL_4P_I1	: in std_logic := '0';
    CAL_4P_I2	: in std_logic := '0';
    CAL_4P_I3	: in std_logic := '0';
    CAL_4P_I4	: in std_logic := '0';
    CAL_4P_I5	: in std_logic := '0';
    CAL_4P_I6	: in std_logic := '0';
    CAL_4P_I7	: in std_logic := '0';
    CAL_4P_I8	: in std_logic := '0';

    CAL_SEL_I1	: in std_logic := '0';
    CAL_SEL_I2	: in std_logic := '0';
    CAL_SEL_I3	: in std_logic := '0';
    CAL_SEL_I4	: in std_logic := '0';

    CAL_E_I	: in std_logic := '0';
    LOCK_E_I	: in std_logic := '0';
    OVS_E_I	: in std_logic := '0';

    TST_I1	: in std_logic := '0';
    TST_I2	: in std_logic := '0';
    TST_I3	: in std_logic := '0';
    TST_I4	: in std_logic := '0';
    TST_I5	: in std_logic := '0';
    TST_I6	: in std_logic := '0';
    TST_I7	: in std_logic := '0';
    TST_I8	: in std_logic := '0';

    CLK_O	: out std_logic := '0';
    LOCK_O	: out std_logic := '0';
    CAL_O	: out std_logic := '0';

    TST_O1	: out std_logic := '0';
    TST_O2	: out std_logic := '0';
    TST_O3	: out std_logic := '0';
    TST_O4	: out std_logic := '0';
    TST_O5	: out std_logic := '0';
    TST_O6	: out std_logic := '0';
    TST_O7	: out std_logic := '0';
    TST_O8	: out std_logic := '0';

    LINK_TX0	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX1	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX2	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX3	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX4	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX5	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX0	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX1	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX2	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX3	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX4	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX5	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');

    CLK_EXT_I	: in std_logic := '0'
);
end component NX_PMA_L;

component NX_CRX_U is
generic (
     cfg_rx_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_on_i                : bit := '0';
     cfg_rx_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_vref_sel_i                  : bit := '0';
     cfg_rx_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_divm_i                      : bit := '0';
     cfg_rx_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_loopback_i                      : bit := '0';
     cfg_rx_pma_clk_pos_i                       : bit := '0';
     cfg_rx_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divm_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divn_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divn_i                      : bit := '0';
     cfg_rx_pcs_debug_en_i                      : bit := '0';
     cfg_rx_pcs_bypass_pma_cdc_i                : bit := '0';
     cfg_rx_pcs_fsm_watchdog_en_i               : bit := '0';
     cfg_rx_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_polarity_i                      : bit := '0';
     cfg_rx_pcs_loopback_i                      : bit := '0';
     cfg_rx_pcs_dscr_bypass_i                   : bit := '0';
     cfg_rx_pcs_8b_dscr_sel_i                   : bit := '0';
     cfg_rx_pcs_replace_bypass_i                : bit := '0';
     cfg_rx_pcs_sync_supported_i                : bit := '0';
     cfg_rx_pcs_buffers_bypass_i                : bit := '0';
     cfg_rx_pcs_buffers_use_cdc_i               : bit := '0';
     cfg_rx_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_only_one_skp_i          : bit := '0';
     cfg_rx_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_dec_bypass_i                    : bit := '0';
     cfg_rx_pcs_align_bypass_i                  : bit := '0';
     cfg_rx_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_en_i                    : bit := '0';
     cfg_rx_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_p_comma_en_i                    : bit := '0';
     cfg_rx_pcs_bypass_usr_cdc_i                : bit := '0';
     cfg_rx_pcs_protocol_size_i                 : bit := '0';
     cfg_rx_gearbox_mode_i                      : bit := '0';
     cfg_rx_gearbox_en_i                        : bit := '0';
     location                     : string := ""
 );
port (
    DSCR_E_I	: in std_logic := '0';
    DEC_E_I	: in std_logic := '0';
    ALIGN_E_I	: in std_logic := '0';
    ALIGN_S_I	: in std_logic := '0';
    REP_E_I	: in std_logic := '0';
    BUF_R_I	: in std_logic := '0';

    OVS_BS_I1	: in std_logic := '0';
    OVS_BS_I2	: in std_logic := '0';

    RST_N_I	: in std_logic := '0';

    PMA_RSTN_I: in  std_logic;
    MEYE_RST_I: in  std_logic;
    PWDN_N_I	: in std_logic := '0';

    DBG_S_I1	: in std_logic := '0';
    DBG_S_I2	: in std_logic := '0';
    DBG_S_I3	: in std_logic := '0';

    DATA_O1	: out std_logic := '0';
    DATA_O2	: out std_logic := '0';
    DATA_O3	: out std_logic := '0';
    DATA_O4	: out std_logic := '0';
    DATA_O5	: out std_logic := '0';
    DATA_O6	: out std_logic := '0';
    DATA_O7	: out std_logic := '0';
    DATA_O8	: out std_logic := '0';
    DATA_O9	: out std_logic := '0';
    DATA_O10	: out std_logic := '0';
    DATA_O11	: out std_logic := '0';
    DATA_O12	: out std_logic := '0';
    DATA_O13	: out std_logic := '0';
    DATA_O14	: out std_logic := '0';
    DATA_O15	: out std_logic := '0';
    DATA_O16	: out std_logic := '0';
    DATA_O17	: out std_logic := '0';
    DATA_O18	: out std_logic := '0';
    DATA_O19	: out std_logic := '0';
    DATA_O20	: out std_logic := '0';
    DATA_O21	: out std_logic := '0';
    DATA_O22	: out std_logic := '0';
    DATA_O23	: out std_logic := '0';
    DATA_O24	: out std_logic := '0';
    DATA_O25	: out std_logic := '0';
    DATA_O26	: out std_logic := '0';
    DATA_O27	: out std_logic := '0';
    DATA_O28	: out std_logic := '0';
    DATA_O29	: out std_logic := '0';
    DATA_O30	: out std_logic := '0';
    DATA_O31	: out std_logic := '0';
    DATA_O32	: out std_logic := '0';
    DATA_O33	: out std_logic := '0';
    DATA_O34	: out std_logic := '0';
    DATA_O35	: out std_logic := '0';
    DATA_O36	: out std_logic := '0';
    DATA_O37	: out std_logic := '0';
    DATA_O38	: out std_logic := '0';
    DATA_O39	: out std_logic := '0';
    DATA_O40	: out std_logic := '0';
    DATA_O41	: out std_logic := '0';
    DATA_O42	: out std_logic := '0';
    DATA_O43	: out std_logic := '0';
    DATA_O44	: out std_logic := '0';
    DATA_O45	: out std_logic := '0';
    DATA_O46	: out std_logic := '0';
    DATA_O47	: out std_logic := '0';
    DATA_O48	: out std_logic := '0';
    DATA_O49	: out std_logic := '0';
    DATA_O50	: out std_logic := '0';
    DATA_O51	: out std_logic := '0';
    DATA_O52	: out std_logic := '0';
    DATA_O53	: out std_logic := '0';
    DATA_O54	: out std_logic := '0';
    DATA_O55	: out std_logic := '0';
    DATA_O56	: out std_logic := '0';
    DATA_O57	: out std_logic := '0';
    DATA_O58	: out std_logic := '0';
    DATA_O59	: out std_logic := '0';
    DATA_O60	: out std_logic := '0';
    DATA_O61	: out std_logic := '0';
    DATA_O62	: out std_logic := '0';
    DATA_O63	: out std_logic := '0';
    DATA_O64	: out std_logic := '0';

    CH_COM_O1	: out std_logic := '0';
    CH_COM_O2	: out std_logic := '0';
    CH_COM_O3	: out std_logic := '0';
    CH_COM_O4	: out std_logic := '0';
    CH_COM_O5	: out std_logic := '0';
    CH_COM_O6	: out std_logic := '0';
    CH_COM_O7	: out std_logic := '0';
    CH_COM_O8	: out std_logic := '0';

    CH_K_O1	: out std_logic := '0';
    CH_K_O2	: out std_logic := '0';
    CH_K_O3	: out std_logic := '0';
    CH_K_O4	: out std_logic := '0';
    CH_K_O5	: out std_logic := '0';
    CH_K_O6	: out std_logic := '0';
    CH_K_O7	: out std_logic := '0';
    CH_K_O8	: out std_logic := '0';

    NIT_O1	: out std_logic := '0';
    NIT_O2	: out std_logic := '0';
    NIT_O3	: out std_logic := '0';
    NIT_O4	: out std_logic := '0';
    NIT_O5	: out std_logic := '0';
    NIT_O6	: out std_logic := '0';
    NIT_O7	: out std_logic := '0';
    NIT_O8	: out std_logic := '0';

    D_ERR_O1	: out std_logic := '0';
    D_ERR_O2	: out std_logic := '0';
    D_ERR_O3	: out std_logic := '0';
    D_ERR_O4	: out std_logic := '0';
    D_ERR_O5	: out std_logic := '0';
    D_ERR_O6	: out std_logic := '0';
    D_ERR_O7	: out std_logic := '0';
    D_ERR_O8	: out std_logic := '0';

    CH_A_O1	: out std_logic := '0';
    CH_A_O2	: out std_logic := '0';
    CH_A_O3	: out std_logic := '0';
    CH_A_O4	: out std_logic := '0';
    CH_A_O5	: out std_logic := '0';
    CH_A_O6	: out std_logic := '0';
    CH_A_O7	: out std_logic := '0';
    CH_A_O8	: out std_logic := '0';

    CH_F_O1	: out std_logic := '0';
    CH_F_O2	: out std_logic := '0';
    CH_F_O3	: out std_logic := '0';
    CH_F_O4	: out std_logic := '0';
    CH_F_O5	: out std_logic := '0';
    CH_F_O6	: out std_logic := '0';
    CH_F_O7	: out std_logic := '0';
    CH_F_O8	: out std_logic := '0';

    ALIGN_O	: out std_logic := '0';
    VREALIGN_O	: out std_logic := '0';
    BUSY_O	: out std_logic := '0';

    TST_O1	: out std_logic := '0';
    TST_O2	: out std_logic := '0';
    TST_O3	: out std_logic := '0';
    TST_O4	: out std_logic := '0';
    TST_O5	: out std_logic := '0';
    TST_O6	: out std_logic := '0';
    TST_O7	: out std_logic := '0';
    TST_O8	: out std_logic := '0';

    LOS_O	: out std_logic := '0';

    LL_FLOCK_O	: out std_logic := '0';
    LL_SLOCK_O	: out std_logic := '0';
    PLL_LOCK_O	: out std_logic := '0';
    PLL_LOCKT_O	: out std_logic := '0';

    LINK	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_CRX_U;

component NX_CTX_U is
generic (
     cfg_tx_pcs_protocol_size_i    : bit := '0';
     cfg_tx_pcs_8b_scr_sel_i       : bit := '0';
     cfg_tx_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
     cfg_tx_pcs_scr_bypass_i       : bit := '0';
     cfg_tx_pcs_sync_supported_i   : bit := '0';
     cfg_tx_pcs_replace_bypass_i   : bit := '0';
     cfg_tx_pcs_enc_bypass_i       : bit := '0';
     cfg_tx_pcs_loopback_i         : bit := '0';
     cfg_tx_pcs_polarity_i         : bit := '0';
     cfg_tx_pcs_esistream_fsm_en_i : bit := '0';
     cfg_tx_pcs_bypass_pma_cdc_i   : bit := '0';
     cfg_tx_pcs_bypass_usr_cdc_i   : bit := '0';
     cfg_tx_pma_clk_pos_i          : bit := '0';
     cfg_tx_pma_loopback_i         : bit := '0';
     cfg_tx_gearbox_en_i           : bit := '0';
     cfg_tx_gearbox_mode_i         : bit := '0';

     location             : string := ""
 );
port (
    ENC_E_I1	: in std_logic := '0';
    ENC_E_I2	: in std_logic := '0';
    ENC_E_I3	: in std_logic := '0';
    ENC_E_I4	: in std_logic := '0';
    ENC_E_I5	: in std_logic := '0';
    ENC_E_I6	: in std_logic := '0';
    ENC_E_I7	: in std_logic := '0';
    ENC_E_I8	: in std_logic := '0';

    CH_K_I1	: in std_logic := '0';
    CH_K_I2	: in std_logic := '0';
    CH_K_I3	: in std_logic := '0';
    CH_K_I4	: in std_logic := '0';
    CH_K_I5	: in std_logic := '0';
    CH_K_I6	: in std_logic := '0';
    CH_K_I7	: in std_logic := '0';
    CH_K_I8	: in std_logic := '0';

    SCR_E_I1	: in std_logic := '0';
    SCR_E_I2	: in std_logic := '0';
    SCR_E_I3	: in std_logic := '0';
    SCR_E_I4	: in std_logic := '0';
    SCR_E_I5	: in std_logic := '0';
    SCR_E_I6	: in std_logic := '0';
    SCR_E_I7	: in std_logic := '0';
    SCR_E_I8	: in std_logic := '0';

    EOMF_I1	: in std_logic := '0';
    EOMF_I2	: in std_logic := '0';
    EOMF_I3	: in std_logic := '0';
    EOMF_I4	: in std_logic := '0';
    EOMF_I5	: in std_logic := '0';
    EOMF_I6	: in std_logic := '0';
    EOMF_I7	: in std_logic := '0';
    EOMF_I8	: in std_logic := '0';

    EOF_I1	: in std_logic := '0';
    EOF_I2	: in std_logic := '0';
    EOF_I3	: in std_logic := '0';
    EOF_I4	: in std_logic := '0';
    EOF_I5	: in std_logic := '0';
    EOF_I6	: in std_logic := '0';
    EOF_I7	: in std_logic := '0';
    EOF_I8	: in std_logic := '0';

    REP_E_I	: in std_logic := '0';
    RST_N_I	: in std_logic := '0';

    DATA_I1	: in std_logic := '0';
    DATA_I2	: in std_logic := '0';
    DATA_I3	: in std_logic := '0';
    DATA_I4	: in std_logic := '0';
    DATA_I5	: in std_logic := '0';
    DATA_I6	: in std_logic := '0';
    DATA_I7	: in std_logic := '0';
    DATA_I8	: in std_logic := '0';
    DATA_I9	: in std_logic := '0';
    DATA_I10	: in std_logic := '0';
    DATA_I11	: in std_logic := '0';
    DATA_I12	: in std_logic := '0';
    DATA_I13	: in std_logic := '0';
    DATA_I14	: in std_logic := '0';
    DATA_I15	: in std_logic := '0';
    DATA_I16	: in std_logic := '0';
    DATA_I17	: in std_logic := '0';
    DATA_I18	: in std_logic := '0';
    DATA_I19	: in std_logic := '0';
    DATA_I20	: in std_logic := '0';
    DATA_I21	: in std_logic := '0';
    DATA_I22	: in std_logic := '0';
    DATA_I23	: in std_logic := '0';
    DATA_I24	: in std_logic := '0';
    DATA_I25	: in std_logic := '0';
    DATA_I26	: in std_logic := '0';
    DATA_I27	: in std_logic := '0';
    DATA_I28	: in std_logic := '0';
    DATA_I29	: in std_logic := '0';
    DATA_I30	: in std_logic := '0';
    DATA_I31	: in std_logic := '0';
    DATA_I32	: in std_logic := '0';
    DATA_I33	: in std_logic := '0';
    DATA_I34	: in std_logic := '0';
    DATA_I35	: in std_logic := '0';
    DATA_I36	: in std_logic := '0';
    DATA_I37	: in std_logic := '0';
    DATA_I38	: in std_logic := '0';
    DATA_I39	: in std_logic := '0';
    DATA_I40	: in std_logic := '0';
    DATA_I41	: in std_logic := '0';
    DATA_I42	: in std_logic := '0';
    DATA_I43	: in std_logic := '0';
    DATA_I44	: in std_logic := '0';
    DATA_I45	: in std_logic := '0';
    DATA_I46	: in std_logic := '0';
    DATA_I47	: in std_logic := '0';
    DATA_I48	: in std_logic := '0';
    DATA_I49	: in std_logic := '0';
    DATA_I50	: in std_logic := '0';
    DATA_I51	: in std_logic := '0';
    DATA_I52	: in std_logic := '0';
    DATA_I53	: in std_logic := '0';
    DATA_I54	: in std_logic := '0';
    DATA_I55	: in std_logic := '0';
    DATA_I56	: in std_logic := '0';
    DATA_I57	: in std_logic := '0';
    DATA_I58	: in std_logic := '0';
    DATA_I59	: in std_logic := '0';
    DATA_I60	: in std_logic := '0';
    DATA_I61	: in std_logic := '0';
    DATA_I62	: in std_logic := '0';
    DATA_I63	: in std_logic := '0';
    DATA_I64	: in std_logic := '0';

    BUSY_O	: out std_logic := '0';
    INV_K_O	: out std_logic := '0';

    PWDN_N_I	: in std_logic := '0';
    CLK_E_I	: in std_logic := '0';

    CLK_O	: out std_logic := '0';

    LINK	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_CTX_U;

component NX_HSSL_U_FULL is
generic (
   -- PMA
   cfg_pll_pma_int_data_len_i            : bit := '0';
   cfg_pll_pma_cpump_i                   : bit_vector( 3 downto 0) := (others => '0');
   cfg_pll_pma_divl_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_divm_i                    : bit := '0';
   cfg_pll_pma_divn_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_lvds_en_i                 : bit := '0';
   cfg_pll_pma_lvds_mux_i                : bit := '0';
   cfg_pll_pma_mux_ckref_i               : bit := '0';
   cfg_pll_pma_gbx_en_i                  : bit := '0';
   cfg_pll_pma_ckref_ext_i               : bit := '0';
   cfg_main_clk_to_fabric_div_mode_i     : bit := '0';
   cfg_main_clk_to_fabric_div_en_i       : bit := '0';
   cfg_main_clk_to_fabric_sel_i          : bit := '0';
   cfg_main_rclk_to_fabric_sel_i         : bit_vector( 1 downto 0) := (others => '0');
   cfg_main_use_only_usr_clock_i         : bit := '0';
   tx_usrclk_use_pcs_clk_2               : bit := '0';
   rx_usrclk_use_pcs_clk_2               : bit := '0';
   cfg_pcs_word_len_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pcs_ovs_en_i                      : bit := '0';
   cfg_pcs_ovs_mode_i                    : bit := '0';
   cfg_pcs_pll_lock_ppm_i                : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_m_eye_i            : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_up_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_dn_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_coarse_ena_i : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_fine_ena_i   : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_step_i       : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_mode_i        : bit_vector( 1 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_locked_i      : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_unlocked_i    : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_1        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_2        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx1_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx2_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx3_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx0_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx1_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx2_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx3_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx0_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_test_mode_i                       : bit_vector( 1 downto 0) := (others => '0');

   --LANE 0
   --TX
   cfg_tx0_pcs_protocol_size_i    : bit := '0';
   cfg_tx0_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx0_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx0_pcs_scr_bypass_i       : bit := '0';
   cfg_tx0_pcs_sync_supported_i   : bit := '0';
   cfg_tx0_pcs_replace_bypass_i   : bit := '0';
   cfg_tx0_pcs_enc_bypass_i       : bit := '0';
   cfg_tx0_pcs_loopback_i         : bit := '0';
   cfg_tx0_pcs_polarity_i         : bit := '0';
   cfg_tx0_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx0_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx0_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx0_pma_clk_pos_i          : bit := '0';
   cfg_tx0_pma_loopback_i         : bit := '0';
   cfg_tx0_gearbox_en_i           : bit := '0';
   cfg_tx0_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx0_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_peak_detect_on_i                : bit := '0';
   cfg_rx0_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx0_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_dco_divm_i                      : bit := '0';
   cfg_rx0_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_loopback_i                      : bit := '0';
   cfg_rx0_pma_clk_pos_i                       : bit := '0';
   cfg_rx0_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divn_i                      : bit := '0';
   cfg_rx0_pcs_debug_en_i                      : bit := '0';
   cfg_rx0_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx0_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx0_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_polarity_i                      : bit := '0';
   cfg_rx0_pcs_loopback_i                      : bit := '0';
   cfg_rx0_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx0_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx0_pcs_replace_bypass_i                : bit := '0';
   cfg_rx0_pcs_sync_supported_i                : bit := '0';
   cfg_rx0_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx0_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx0_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx0_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx0_pcs_align_bypass_i                  : bit := '0';
   cfg_rx0_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx0_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx0_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx0_pcs_protocol_size_i                 : bit := '0';
   cfg_rx0_gearbox_mode_i                      : bit := '0';
   cfg_rx0_gearbox_en_i                        : bit := '0';

   --LANE 1
   --TX
   cfg_tx1_pcs_protocol_size_i    : bit := '0';
   cfg_tx1_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx1_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx1_pcs_scr_bypass_i       : bit := '0';
   cfg_tx1_pcs_sync_supported_i   : bit := '0';
   cfg_tx1_pcs_replace_bypass_i   : bit := '0';
   cfg_tx1_pcs_enc_bypass_i       : bit := '0';
   cfg_tx1_pcs_loopback_i         : bit := '0';
   cfg_tx1_pcs_polarity_i         : bit := '0';
   cfg_tx1_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx1_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx1_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx1_pma_clk_pos_i          : bit := '0';
   cfg_tx1_pma_loopback_i         : bit := '0';
   cfg_tx1_gearbox_en_i           : bit := '0';
   cfg_tx1_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx1_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_peak_detect_on_i                : bit := '0';
   cfg_rx1_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx1_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_dco_divm_i                      : bit := '0';
   cfg_rx1_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_loopback_i                      : bit := '0';
   cfg_rx1_pma_clk_pos_i                       : bit := '0';
   cfg_rx1_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divn_i                      : bit := '0';
   cfg_rx1_pcs_debug_en_i                      : bit := '0';
   cfg_rx1_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx1_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx1_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_polarity_i                      : bit := '0';
   cfg_rx1_pcs_loopback_i                      : bit := '0';
   cfg_rx1_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx1_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx1_pcs_replace_bypass_i                : bit := '0';
   cfg_rx1_pcs_sync_supported_i                : bit := '0';
   cfg_rx1_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx1_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx1_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx1_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx1_pcs_align_bypass_i                  : bit := '0';
   cfg_rx1_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx1_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx1_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx1_pcs_protocol_size_i                 : bit := '0';
   cfg_rx1_gearbox_mode_i                      : bit := '0';
   cfg_rx1_gearbox_en_i                        : bit := '0';

   --LANE 2
   --TX
   cfg_tx2_pcs_protocol_size_i    : bit := '0';
   cfg_tx2_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx2_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx2_pcs_scr_bypass_i       : bit := '0';
   cfg_tx2_pcs_sync_supported_i   : bit := '0';
   cfg_tx2_pcs_replace_bypass_i   : bit := '0';
   cfg_tx2_pcs_enc_bypass_i       : bit := '0';
   cfg_tx2_pcs_loopback_i         : bit := '0';
   cfg_tx2_pcs_polarity_i         : bit := '0';
   cfg_tx2_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx2_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx2_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx2_pma_clk_pos_i          : bit := '0';
   cfg_tx2_pma_loopback_i         : bit := '0';
   cfg_tx2_gearbox_en_i           : bit := '0';
   cfg_tx2_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx2_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_peak_detect_on_i                : bit := '0';
   cfg_rx2_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx2_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_dco_divm_i                      : bit := '0';
   cfg_rx2_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_loopback_i                      : bit := '0';
   cfg_rx2_pma_clk_pos_i                       : bit := '0';
   cfg_rx2_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divn_i                      : bit := '0';
   cfg_rx2_pcs_debug_en_i                      : bit := '0';
   cfg_rx2_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx2_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx2_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_polarity_i                      : bit := '0';
   cfg_rx2_pcs_loopback_i                      : bit := '0';
   cfg_rx2_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx2_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx2_pcs_replace_bypass_i                : bit := '0';
   cfg_rx2_pcs_sync_supported_i                : bit := '0';
   cfg_rx2_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx2_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx2_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx2_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx2_pcs_align_bypass_i                  : bit := '0';
   cfg_rx2_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx2_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx2_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx2_pcs_protocol_size_i                 : bit := '0';
   cfg_rx2_gearbox_mode_i                      : bit := '0';
   cfg_rx2_gearbox_en_i                        : bit := '0';

   --LANE 3
   --TX
   cfg_tx3_pcs_protocol_size_i    : bit := '0';
   cfg_tx3_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx3_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx3_pcs_scr_bypass_i       : bit := '0';
   cfg_tx3_pcs_sync_supported_i   : bit := '0';
   cfg_tx3_pcs_replace_bypass_i   : bit := '0';
   cfg_tx3_pcs_enc_bypass_i       : bit := '0';
   cfg_tx3_pcs_loopback_i         : bit := '0';
   cfg_tx3_pcs_polarity_i         : bit := '0';
   cfg_tx3_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx3_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx3_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx3_pma_clk_pos_i          : bit := '0';
   cfg_tx3_pma_loopback_i         : bit := '0';
   cfg_tx3_gearbox_en_i           : bit := '0';
   cfg_tx3_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx3_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_peak_detect_on_i                : bit := '0';
   cfg_rx3_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx3_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_dco_divm_i                      : bit := '0';
   cfg_rx3_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_loopback_i                      : bit := '0';
   cfg_rx3_pma_clk_pos_i                       : bit := '0';
   cfg_rx3_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divn_i                      : bit := '0';
   cfg_rx3_pcs_debug_en_i                      : bit := '0';
   cfg_rx3_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx3_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx3_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_polarity_i                      : bit := '0';
   cfg_rx3_pcs_loopback_i                      : bit := '0';
   cfg_rx3_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx3_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx3_pcs_replace_bypass_i                : bit := '0';
   cfg_rx3_pcs_sync_supported_i                : bit := '0';
   cfg_rx3_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx3_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx3_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx3_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx3_pcs_align_bypass_i                  : bit := '0';
   cfg_rx3_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx3_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx3_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx3_pcs_protocol_size_i                 : bit := '0';
   cfg_rx3_gearbox_mode_i                      : bit := '0';
   cfg_rx3_gearbox_en_i                        : bit := '0';

   location   : string := ""
 );
port (
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ MAIN ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- PMA
    hssl_clk_user_tx_i	: in std_logic := '0';
    hssl_clk_user_rx_i	: in std_logic := '0';
    hssl_clk_ref_i	: in std_logic := '0';
    hssl_clock_o	: out std_logic := '0';
    hssl_rclock_o	: out std_logic := '0';
    usr_dyn_cfg_en_i	: in std_logic := '0';
    usr_dyn_cfg_lane_cs_n_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_dyn_cfg_calibration_cs_n_i	: in std_logic := '0';
    usr_dyn_cfg_we_n_i	: in std_logic := '0';
    usr_dyn_cfg_addr_i	: in std_logic_vector(3 downto 0) := (others => '0');
    usr_dyn_cfg_wdata_sel_i	: in std_logic := '0';
    usr_dyn_cfg_wdata_i	: in std_logic_vector(11 downto 0) := (others => '0');
    usr_pll_pma_rst_n_i	: in std_logic := '0';
    usr_pll_pma_pwr_down_n_i	: in std_logic := '0';
    usr_main_rst_n_i	: in std_logic := '0';
    usr_pll_lock_o	: out std_logic := '0';
    usr_pll_pma_lock_analog_o	: out std_logic := '0';
    usr_pll_ckfb_lock_o	: out std_logic := '0';
    usr_calibrate_pma_out_o	: out std_logic := '0';
    usr_main_async_debug_lane_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_main_async_debug_ack_i	: in std_logic := '0';
    usr_main_async_debug_req_o	: out std_logic := '0';
    usr_main_rx_pma_ll_out_o	: out std_logic_vector(19 downto 0) := (others => '0');
    scan_en_i	: in std_logic := '0';
    scan_in_i	: in std_logic_vector(7 downto 0) := (others => '0');
    scan_out_o	: out std_logic_vector(7 downto 0) := (others => '0');


   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 0 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
    usr_tx0_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx0_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx0_rst_n_i	: in std_logic := '0';
    usr_tx0_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx0_busy_o	: out std_logic := '0';
    usr_tx0_ctrl_invalid_k_o	: out std_logic := '0';
    usr_tx0_ctrl_driver_pwrdwn_n_i	: in std_logic := '0';
    usr_tx0_pma_clk_en_i	: in std_logic := '0';
    usr_tx0_pma_tx_clk_o	: out std_logic := '0';

    -- RX - Fabric Interface
    usr_rx0_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx0_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx0_ctrl_align_en_i	: in std_logic := '0';
    usr_rx0_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx0_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx0_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx0_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx0_rst_n_i	: in std_logic := '0';
    usr_rx0_pma_rst_n_i	: in std_logic := '0';
    usr_rx0_pma_m_eye_rst_i	: in std_logic := '0';
    usr_rx0_pma_pwr_down_n_i	: in std_logic := '0';
    usr_rx0_ctrl_debug_sel_i	: in std_logic_vector(2 downto 0) := (others => '0');
    usr_rx0_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx0_ctrl_valid_realign_o	: out std_logic := '0';
    usr_rx0_busy_o	: out std_logic := '0';
    usr_rx0_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx0_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx0_pma_ll_fast_locked_o	: out std_logic := '0';
    usr_rx0_pma_ll_slow_locked_o	: out std_logic := '0';
    usr_rx0_pma_pll_lock_o	: out std_logic := '0';
    usr_rx0_pma_pll_lock_track_o	: out std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 1 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
    usr_tx1_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx1_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx1_rst_n_i	: in std_logic := '0';
    usr_tx1_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx1_busy_o	: out std_logic := '0';
    usr_tx1_ctrl_invalid_k_o	: out std_logic := '0';
    usr_tx1_ctrl_driver_pwrdwn_n_i	: in std_logic := '0';
    usr_tx1_pma_clk_en_i	: in std_logic := '0';
    usr_tx1_pma_tx_clk_o	: out std_logic := '0';

    -- RX - Fabric Interface
    usr_rx1_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx1_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx1_ctrl_align_en_i	: in std_logic := '0';
    usr_rx1_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx1_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx1_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx1_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx1_rst_n_i	: in std_logic := '0';
    usr_rx1_pma_rst_n_i	: in std_logic := '0';
    usr_rx1_pma_m_eye_rst_i	: in std_logic := '0';
    usr_rx1_pma_pwr_down_n_i	: in std_logic := '0';
    usr_rx1_ctrl_debug_sel_i	: in std_logic_vector(2 downto 0) := (others => '0');
    usr_rx1_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx1_ctrl_valid_realign_o	: out std_logic := '0';
    usr_rx1_busy_o	: out std_logic := '0';
    usr_rx1_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx1_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx1_pma_ll_fast_locked_o	: out std_logic := '0';
    usr_rx1_pma_ll_slow_locked_o	: out std_logic := '0';
    usr_rx1_pma_pll_lock_o	: out std_logic := '0';
    usr_rx1_pma_pll_lock_track_o	: out std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 2 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
    usr_tx2_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx2_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx2_rst_n_i	: in std_logic := '0';
    usr_tx2_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx2_busy_o	: out std_logic := '0';
    usr_tx2_ctrl_invalid_k_o	: out std_logic := '0';
    usr_tx2_ctrl_driver_pwrdwn_n_i	: in std_logic := '0';
    usr_tx2_pma_clk_en_i	: in std_logic := '0';
    usr_tx2_pma_tx_clk_o	: out std_logic := '0';

   -- RX - Fabric Interface
    usr_rx2_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx2_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx2_ctrl_align_en_i	: in std_logic := '0';
    usr_rx2_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx2_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx2_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx2_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx2_rst_n_i	: in std_logic := '0';
    usr_rx2_pma_rst_n_i	: in std_logic := '0';
    usr_rx2_pma_m_eye_rst_i	: in std_logic := '0';
    usr_rx2_pma_pwr_down_n_i	: in std_logic := '0';
    usr_rx2_ctrl_debug_sel_i	: in std_logic_vector(2 downto 0) := (others => '0');
    usr_rx2_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx2_ctrl_valid_realign_o	: out std_logic := '0';
    usr_rx2_busy_o	: out std_logic := '0';
    usr_rx2_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx2_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx2_pma_ll_fast_locked_o	: out std_logic := '0';
    usr_rx2_pma_ll_slow_locked_o	: out std_logic := '0';
    usr_rx2_pma_pll_lock_o	: out std_logic := '0';
    usr_rx2_pma_pll_lock_track_o	: out std_logic := '0';

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 3 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
    usr_tx3_ctrl_enc_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_char_is_k_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_scr_en_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_end_of_multiframe_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_end_of_frame_i	: in std_logic_vector(7 downto 0) := (others => '0');
    usr_tx3_ctrl_replace_en_i	: in std_logic := '0';
    usr_tx3_rst_n_i	: in std_logic := '0';
    usr_tx3_data_i	: in std_logic_vector(63 downto 0) := (others => '0');
    usr_tx3_busy_o	: out std_logic := '0';
    usr_tx3_ctrl_invalid_k_o	: out std_logic := '0';
    usr_tx3_ctrl_driver_pwrdwn_n_i	: in std_logic := '0';
    usr_tx3_pma_clk_en_i	: in std_logic := '0';
    usr_tx3_pma_tx_clk_o	: out std_logic := '0';

   -- RX - Fabric Interface
    usr_rx3_ctrl_dscr_en_i	: in std_logic := '0';
    usr_rx3_ctrl_dec_en_i	: in std_logic := '0';
    usr_rx3_ctrl_align_en_i	: in std_logic := '0';
    usr_rx3_ctrl_align_sync_i	: in std_logic := '0';
    usr_rx3_ctrl_replace_en_i	: in std_logic := '0';
    usr_rx3_ctrl_el_buff_rst_i	: in std_logic := '0';
    usr_rx3_ctrl_ovs_bit_sel_i	: in std_logic_vector(1 downto 0) := (others => '0');
    usr_rx3_rst_n_i	: in std_logic := '0';
    usr_rx3_pma_rst_n_i	: in std_logic := '0';
    usr_rx3_pma_m_eye_rst_i	: in std_logic := '0';
    usr_rx3_pma_pwr_down_n_i	: in std_logic := '0';
    usr_rx3_ctrl_debug_sel_i	: in std_logic_vector(2 downto 0) := (others => '0');
    usr_rx3_data_o	: out std_logic_vector(63 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_comma_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_k_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_not_in_table_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_disp_err_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_a_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_f_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_ctrl_char_is_aligned_o	: out std_logic := '0';
    usr_rx3_ctrl_valid_realign_o	: out std_logic := '0';
    usr_rx3_busy_o	: out std_logic := '0';
    usr_rx3_test_o	: out std_logic_vector(7 downto 0) := (others => '0');
    usr_rx3_pma_loss_of_signal_o	: out std_logic := '0';
    usr_rx3_pma_ll_fast_locked_o	: out std_logic := '0';
    usr_rx3_pma_ll_slow_locked_o	: out std_logic := '0';
    usr_rx3_pma_pll_lock_o	: out std_logic := '0';
    usr_rx3_pma_pll_lock_track_o	: out std_logic := '0'
);
end component NX_HSSL_U_FULL;

component NX_PMA_U is
generic (
   cfg_pll_pma_int_data_len_i            : bit := '0';
   cfg_pll_pma_cpump_i                   : bit_vector( 3 downto 0) := (others => '0');
   cfg_pll_pma_divl_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_divm_i                    : bit := '0';
   cfg_pll_pma_divn_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_lvds_en_i                 : bit := '0';
   cfg_pll_pma_lvds_mux_i                : bit := '0';
   cfg_pll_pma_mux_ckref_i               : bit := '0';
   cfg_pll_pma_gbx_en_i                  : bit := '0';
   cfg_pll_pma_ckref_ext_i               : bit := '0';
   cfg_main_clk_to_fabric_div_mode_i     : bit := '0';
   cfg_main_clk_to_fabric_div_en_i       : bit := '0';
   cfg_main_clk_to_fabric_sel_i          : bit := '0';
   cfg_main_rclk_to_fabric_sel_i         : bit_vector( 1 downto 0) := (others => '0');
   cfg_main_use_only_usr_clock_i         : bit := '0';
   tx_usrclk_use_pcs_clk_2               : bit := '0';
   rx_usrclk_use_pcs_clk_2               : bit := '0';
   cfg_pcs_word_len_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pcs_ovs_en_i                      : bit := '0';
   cfg_pcs_ovs_mode_i                    : bit := '0';
   cfg_pcs_pll_lock_ppm_i                : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_m_eye_i            : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_up_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_dn_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_coarse_ena_i : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_fine_ena_i   : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_step_i       : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_mode_i        : bit_vector( 1 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_locked_i      : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_unlocked_i    : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_1        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_2        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx1_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx2_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx3_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx0_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx1_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx2_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx3_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx0_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_test_mode_i                       : bit_vector( 1 downto 0) := (others => '0');

   location                    : string := ""
);
port (
    CLK_TX_I	: in std_logic := '0';
    CLK_RX_I	: in std_logic := '0';
    CLK_REF_I	: in std_logic := '0';

    DC_E_I	: in std_logic := '0';
    DC_LCSN_I1	: in std_logic := '0';
    DC_LCSN_I2	: in std_logic := '0';
    DC_LCSN_I3	: in std_logic := '0';
    DC_LCSN_I4	: in std_logic := '0';

    DC_CCSN_I	: in std_logic := '0';
    DC_WE_N_I	: in std_logic := '0';

    DC_ADD_I1	: in std_logic := '0';
    DC_ADD_I2	: in std_logic := '0';
    DC_ADD_I3	: in std_logic := '0';
    DC_ADD_I4	: in std_logic := '0';
    DC_WDATAS_I	: in std_logic := '0';
    DC_WDATA_I1	: in std_logic := '0';
    DC_WDATA_I2	: in std_logic := '0';
    DC_WDATA_I3	: in std_logic := '0';
    DC_WDATA_I4	: in std_logic := '0';
    DC_WDATA_I5	: in std_logic := '0';
    DC_WDATA_I6	: in std_logic := '0';
    DC_WDATA_I7	: in std_logic := '0';
    DC_WDATA_I8	: in std_logic := '0';
    DC_WDATA_I9	: in std_logic := '0';
    DC_WDATA_I10	: in std_logic := '0';
    DC_WDATA_I11	: in std_logic := '0';
    DC_WDATA_I12	: in std_logic := '0';

    PLL_RN_I	: in std_logic := '0';
    PWDN_N_I	: in std_logic := '0';
    RST_N_I	: in std_logic := '0';

    DBG_S_I1	: in std_logic := '0';
    DBG_S_I2	: in std_logic := '0';
    DBG_A_I	: in std_logic := '0';

    SE_I	: in std_logic := '0';

    SCAN_I1	: in std_logic := '0';
    SCAN_I2	: in std_logic := '0';
    SCAN_I3	: in std_logic := '0';
    SCAN_I4	: in std_logic := '0';
    SCAN_I5	: in std_logic := '0';
    SCAN_I6	: in std_logic := '0';
    SCAN_I7	: in std_logic := '0';
    SCAN_I8	: in std_logic := '0';

    CLK_O	: out std_logic := '0';
    CLK_RX_O	: out std_logic := '0';
    LOCK_O	: out std_logic := '0';
    LOCKA_O	: out std_logic := '0';
    FB_LOCK_O	: out std_logic := '0';
    CAL_OUT_O	: out std_logic := '0';
    DBG_R_O	: out std_logic := '0';

    LL_O1	: out std_logic := '0';
    LL_O2	: out std_logic := '0';
    LL_O3	: out std_logic := '0';
    LL_O4	: out std_logic := '0';
    LL_O5	: out std_logic := '0';
    LL_O6	: out std_logic := '0';
    LL_O7	: out std_logic := '0';
    LL_O8	: out std_logic := '0';
    LL_O9	: out std_logic := '0';
    LL_O10	: out std_logic := '0';
    LL_O11	: out std_logic := '0';
    LL_O12	: out std_logic := '0';
    LL_O13	: out std_logic := '0';
    LL_O14	: out std_logic := '0';
    LL_O15	: out std_logic := '0';
    LL_O16	: out std_logic := '0';
    LL_O17	: out std_logic := '0';
    LL_O18	: out std_logic := '0';
    LL_O19	: out std_logic := '0';
    LL_O20	: out std_logic := '0';


    SCAN_O1	: out std_logic := '0';
    SCAN_O2	: out std_logic := '0';
    SCAN_O3	: out std_logic := '0';
    SCAN_O4	: out std_logic := '0';
    SCAN_O5	: out std_logic := '0';
    SCAN_O6	: out std_logic := '0';
    SCAN_O7	: out std_logic := '0';
    SCAN_O8	: out std_logic := '0';


    LINK_TX0	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX1	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX2	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_TX3	: inout std_logic_vector(CTX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX0	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX1	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX2	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0');
    LINK_RX3	: inout std_logic_vector(CRX_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_PMA_U;

component NX_IOM_L is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk1 : bit := '0';
--  latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk2 : bit := '0';
--  latency2     : bit := '0';
--  sel_clk_out2 : bit_vector(1 downto 0) := "00";
--  sel_clk_out3 : bit_vector(1 downto 0) := "00";
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_io_cal  : bit := '0';
    pads_dict    : string := "";
    pads_path    : string := ""
);
port (
    RTCK1	: in std_logic := '0';
    RRCK1	: in std_logic := '0';
    WTCK1	: in std_logic := '0';
    WRCK1	: in std_logic := '0';
    RTCK2	: in std_logic := '0';
    RRCK2	: in std_logic := '0';
    WTCK2	: in std_logic := '0';
    WRCK2	: in std_logic := '0';
    CTCK	: in std_logic := '0';
    CCK	: in std_logic := '0';
    DCK	: in std_logic := '0';

    C1TW	: in std_logic := '0';
    C1TS	: in std_logic := '0';
    C1RW1	: in std_logic := '0';
    C1RW2	: in std_logic := '0';
    C1RW3	: in std_logic := '0';
    C1RNE	: in std_logic := '0';
    C1RS	: in std_logic := '0';
    C2TW	: in std_logic := '0';
    C2TS	: in std_logic := '0';
    C2RW1	: in std_logic := '0';
    C2RW2	: in std_logic := '0';
    C2RW3	: in std_logic := '0';
    C2RNE	: in std_logic := '0';
    C2RS	: in std_logic := '0';
    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';
    DC	: in std_logic := '0';
    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';
    DRA5	: in std_logic := '0';
    DRA6	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DOS	: in std_logic := '0';
    DOG	: in std_logic := '0';
    DIS	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DPAS	: in std_logic := '0';
    DPAG	: in std_logic := '0';
    DQSS	: in std_logic := '0';
    DQSG	: in std_logic := '0';
    DS1	: in std_logic := '0';
    DS2	: in std_logic := '0';
    CAD1	: in std_logic := '0';
    CAD2	: in std_logic := '0';
    CAD3	: in std_logic := '0';
    CAD4	: in std_logic := '0';
    CAD5	: in std_logic := '0';
    CAD6	: in std_logic := '0';
    CAP1	: in std_logic := '0';
    CAP2	: in std_logic := '0';
    CAP3	: in std_logic := '0';
    CAP4	: in std_logic := '0';
    CAN1	: in std_logic := '0';
    CAN2	: in std_logic := '0';
    CAN3	: in std_logic := '0';
    CAN4	: in std_logic := '0';
    CAT1	: in std_logic := '0';
    CAT2	: in std_logic := '0';
    CAT3	: in std_logic := '0';
    CAT4	: in std_logic := '0';

    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';

    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    C1RED	: out std_logic := '0';
    C2RED	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';
    CAL	: out std_logic := '0';

    P1CI1	: in std_logic := '0';
    P1CL	: in std_logic := '0';
    P1CR	: in std_logic := '0';
    P1CO	: out std_logic := '0';
    P1CTI	: in std_logic := '0';
    P1CTO	: out std_logic := '0';
    P1EI1	: in std_logic := '0';
    P1EI2	: in std_logic := '0';
    P1EI3	: in std_logic := '0';
    P1EI4	: in std_logic := '0';
    P1EI5	: in std_logic := '0';
    P1EL	: in std_logic := '0';
    P1ER	: in std_logic := '0';
    P1EO	: out std_logic := '0';
    P1RI	: in std_logic := '0';
    P1RL	: in std_logic := '0';
    P1RR	: in std_logic := '0';
    P1RO1	: out std_logic := '0';
    P1RO2	: out std_logic := '0';
    P1RO3	: out std_logic := '0';
    P1RO4	: out std_logic := '0';
    P1RO5	: out std_logic := '0';

    P2CI1	: in std_logic := '0';
    P2CL	: in std_logic := '0';
    P2CR	: in std_logic := '0';
    P2CO	: out std_logic := '0';
    P2CTI	: in std_logic := '0';
    P2CTO	: out std_logic := '0';
    P2EI1	: in std_logic := '0';
    P2EI2	: in std_logic := '0';
    P2EI3	: in std_logic := '0';
    P2EI4	: in std_logic := '0';
    P2EI5	: in std_logic := '0';
    P2EL	: in std_logic := '0';
    P2ER	: in std_logic := '0';
    P2EO	: out std_logic := '0';
    P2RI	: in std_logic := '0';
    P2RL	: in std_logic := '0';
    P2RR	: in std_logic := '0';
    P2RO1	: out std_logic := '0';
    P2RO2	: out std_logic := '0';
    P2RO3	: out std_logic := '0';
    P2RO4	: out std_logic := '0';
    P2RO5	: out std_logic := '0';

    P3CI1	: in std_logic := '0';
    P3CL	: in std_logic := '0';
    P3CR	: in std_logic := '0';
    P3CO	: out std_logic := '0';
    P3CTI	: in std_logic := '0';
    P3CTO	: out std_logic := '0';
    P3EI1	: in std_logic := '0';
    P3EI2	: in std_logic := '0';
    P3EI3	: in std_logic := '0';
    P3EI4	: in std_logic := '0';
    P3EI5	: in std_logic := '0';
    P3EL	: in std_logic := '0';
    P3ER	: in std_logic := '0';
    P3EO	: out std_logic := '0';
    P3RI	: in std_logic := '0';
    P3RL	: in std_logic := '0';
    P3RR	: in std_logic := '0';
    P3RO1	: out std_logic := '0';
    P3RO2	: out std_logic := '0';
    P3RO3	: out std_logic := '0';
    P3RO4	: out std_logic := '0';
    P3RO5	: out std_logic := '0';

    P4CI1	: in std_logic := '0';
    P4CL	: in std_logic := '0';
    P4CR	: in std_logic := '0';
    P4CO	: out std_logic := '0';
    P4CTI	: in std_logic := '0';
    P4CTO	: out std_logic := '0';
    P4EI1	: in std_logic := '0';
    P4EI2	: in std_logic := '0';
    P4EI3	: in std_logic := '0';
    P4EI4	: in std_logic := '0';
    P4EI5	: in std_logic := '0';
    P4EL	: in std_logic := '0';
    P4ER	: in std_logic := '0';
    P4EO	: out std_logic := '0';
    P4RI	: in std_logic := '0';
    P4RL	: in std_logic := '0';
    P4RR	: in std_logic := '0';
    P4RO1	: out std_logic := '0';
    P4RO2	: out std_logic := '0';
    P4RO3	: out std_logic := '0';
    P4RO4	: out std_logic := '0';
    P4RO5	: out std_logic := '0';

    P5CI1	: in std_logic := '0';
    P5CI2	: in std_logic := '0';
    P5CI3	: in std_logic := '0';
    P5CI4	: in std_logic := '0';
    P5CI5	: in std_logic := '0';
    P5CL	: in std_logic := '0';
    P5CR	: in std_logic := '0';
    P5CO	: out std_logic := '0';
    P5CTI	: in std_logic := '0';
    P5CTO	: out std_logic := '0';
    P5EI1	: in std_logic := '0';
    P5EI2	: in std_logic := '0';
    P5EI3	: in std_logic := '0';
    P5EI4	: in std_logic := '0';
    P5EI5	: in std_logic := '0';
    P5EL	: in std_logic := '0';
    P5ER	: in std_logic := '0';
    P5EO	: out std_logic := '0';
    P5RI	: in std_logic := '0';
    P5RL	: in std_logic := '0';
    P5RR	: in std_logic := '0';
    P5RO1	: out std_logic := '0';
    P5RO2	: out std_logic := '0';
    P5RO3	: out std_logic := '0';
    P5RO4	: out std_logic := '0';
    P5RO5	: out std_logic := '0';

    P6CI1	: in std_logic := '0';
    P6CL	: in std_logic := '0';
    P6CR	: in std_logic := '0';
    P6CO	: out std_logic := '0';
    P6CTI	: in std_logic := '0';
    P6CTO	: out std_logic := '0';
    P6EI1	: in std_logic := '0';
    P6EI2	: in std_logic := '0';
    P6EI3	: in std_logic := '0';
    P6EI4	: in std_logic := '0';
    P6EI5	: in std_logic := '0';
    P6EL	: in std_logic := '0';
    P6ER	: in std_logic := '0';
    P6EO	: out std_logic := '0';
    P6RI	: in std_logic := '0';
    P6RL	: in std_logic := '0';
    P6RR	: in std_logic := '0';
    P6RO1	: out std_logic := '0';
    P6RO2	: out std_logic := '0';
    P6RO3	: out std_logic := '0';
    P6RO4	: out std_logic := '0';
    P6RO5	: out std_logic := '0';

    P7CI1	: in std_logic := '0';
    P7CL	: in std_logic := '0';
    P7CR	: in std_logic := '0';
    P7CO	: out std_logic := '0';
    P7CTI	: in std_logic := '0';
    P7CTO	: out std_logic := '0';
    P7EI1	: in std_logic := '0';
    P7EI2	: in std_logic := '0';
    P7EI3	: in std_logic := '0';
    P7EI4	: in std_logic := '0';
    P7EI5	: in std_logic := '0';
    P7EL	: in std_logic := '0';
    P7ER	: in std_logic := '0';
    P7EO	: out std_logic := '0';
    P7RI	: in std_logic := '0';
    P7RL	: in std_logic := '0';
    P7RR	: in std_logic := '0';
    P7RO1	: out std_logic := '0';
    P7RO2	: out std_logic := '0';
    P7RO3	: out std_logic := '0';
    P7RO4	: out std_logic := '0';
    P7RO5	: out std_logic := '0';

    P8CI1	: in std_logic := '0';
    P8CL	: in std_logic := '0';
    P8CR	: in std_logic := '0';
    P8CO	: out std_logic := '0';
    P8CTI	: in std_logic := '0';
    P8CTO	: out std_logic := '0';
    P8EI1	: in std_logic := '0';
    P8EI2	: in std_logic := '0';
    P8EI3	: in std_logic := '0';
    P8EI4	: in std_logic := '0';
    P8EI5	: in std_logic := '0';
    P8EL	: in std_logic := '0';
    P8ER	: in std_logic := '0';
    P8EO	: out std_logic := '0';
    P8RI	: in std_logic := '0';
    P8RL	: in std_logic := '0';
    P8RR	: in std_logic := '0';
    P8RO1	: out std_logic := '0';
    P8RO2	: out std_logic := '0';
    P8RO3	: out std_logic := '0';
    P8RO4	: out std_logic := '0';
    P8RO5	: out std_logic := '0';

    P9CI1	: in std_logic := '0';
    P9CL	: in std_logic := '0';
    P9CR	: in std_logic := '0';
    P9CO	: out std_logic := '0';
    P9CTI	: in std_logic := '0';
    P9CTO	: out std_logic := '0';
    P9EI1	: in std_logic := '0';
    P9EI2	: in std_logic := '0';
    P9EI3	: in std_logic := '0';
    P9EI4	: in std_logic := '0';
    P9EI5	: in std_logic := '0';
    P9EL	: in std_logic := '0';
    P9ER	: in std_logic := '0';
    P9EO	: out std_logic := '0';
    P9RI	: in std_logic := '0';
    P9RL	: in std_logic := '0';
    P9RR	: in std_logic := '0';
    P9RO1	: out std_logic := '0';
    P9RO2	: out std_logic := '0';
    P9RO3	: out std_logic := '0';
    P9RO4	: out std_logic := '0';
    P9RO5	: out std_logic := '0';

    P10CI1	: in std_logic := '0';
    P10CL	: in std_logic := '0';
    P10CR	: in std_logic := '0';
    P10CO	: out std_logic := '0';
    P10CTI	: in std_logic := '0';
    P10CTO	: out std_logic := '0';
    P10EI1	: in std_logic := '0';
    P10EI2	: in std_logic := '0';
    P10EI3	: in std_logic := '0';
    P10EI4	: in std_logic := '0';
    P10EI5	: in std_logic := '0';
    P10EL	: in std_logic := '0';
    P10ER	: in std_logic := '0';
    P10EO	: out std_logic := '0';
    P10RI	: in std_logic := '0';
    P10RL	: in std_logic := '0';
    P10RR	: in std_logic := '0';
    P10RO1	: out std_logic := '0';
    P10RO2	: out std_logic := '0';
    P10RO3	: out std_logic := '0';
    P10RO4	: out std_logic := '0';
    P10RO5	: out std_logic := '0';

    P11CI1	: in std_logic := '0';
    P11CL	: in std_logic := '0';
    P11CR	: in std_logic := '0';
    P11CO	: out std_logic := '0';
    P11CTI	: in std_logic := '0';
    P11CTO	: out std_logic := '0';
    P11EI1	: in std_logic := '0';
    P11EI2	: in std_logic := '0';
    P11EI3	: in std_logic := '0';
    P11EI4	: in std_logic := '0';
    P11EI5	: in std_logic := '0';
    P11EL	: in std_logic := '0';
    P11ER	: in std_logic := '0';
    P11EO	: out std_logic := '0';
    P11RI	: in std_logic := '0';
    P11RL	: in std_logic := '0';
    P11RR	: in std_logic := '0';
    P11RO1	: out std_logic := '0';
    P11RO2	: out std_logic := '0';
    P11RO3	: out std_logic := '0';
    P11RO4	: out std_logic := '0';
    P11RO5	: out std_logic := '0';

    P12CI1	: in std_logic := '0';
    P12CL	: in std_logic := '0';
    P12CR	: in std_logic := '0';
    P12CO	: out std_logic := '0';
    P12CTI	: in std_logic := '0';
    P12CTO	: out std_logic := '0';
    P12EI1	: in std_logic := '0';
    P12EI2	: in std_logic := '0';
    P12EI3	: in std_logic := '0';
    P12EI4	: in std_logic := '0';
    P12EI5	: in std_logic := '0';
    P12EL	: in std_logic := '0';
    P12ER	: in std_logic := '0';
    P12EO	: out std_logic := '0';
    P12RI	: in std_logic := '0';
    P12RL	: in std_logic := '0';
    P12RR	: in std_logic := '0';
    P12RO1	: out std_logic := '0';
    P12RO2	: out std_logic := '0';
    P12RO3	: out std_logic := '0';
    P12RO4	: out std_logic := '0';
    P12RO5	: out std_logic := '0';

    P13CI1	: in std_logic := '0';
    P13CL	: in std_logic := '0';
    P13CR	: in std_logic := '0';
    P13CO	: out std_logic := '0';
    P13CTI	: in std_logic := '0';
    P13CTO	: out std_logic := '0';
    P13EI1	: in std_logic := '0';
    P13EI2	: in std_logic := '0';
    P13EI3	: in std_logic := '0';
    P13EI4	: in std_logic := '0';
    P13EI5	: in std_logic := '0';
    P13EL	: in std_logic := '0';
    P13ER	: in std_logic := '0';
    P13EO	: out std_logic := '0';
    P13RI	: in std_logic := '0';
    P13RL	: in std_logic := '0';
    P13RR	: in std_logic := '0';
    P13RO1	: out std_logic := '0';
    P13RO2	: out std_logic := '0';
    P13RO3	: out std_logic := '0';
    P13RO4	: out std_logic := '0';
    P13RO5	: out std_logic := '0';

    P14CI1	: in std_logic := '0';
    P14CL	: in std_logic := '0';
    P14CR	: in std_logic := '0';
    P14CO	: out std_logic := '0';
    P14CTI	: in std_logic := '0';
    P14CTO	: out std_logic := '0';
    P14EI1	: in std_logic := '0';
    P14EI2	: in std_logic := '0';
    P14EI3	: in std_logic := '0';
    P14EI4	: in std_logic := '0';
    P14EI5	: in std_logic := '0';
    P14EL	: in std_logic := '0';
    P14ER	: in std_logic := '0';
    P14EO	: out std_logic := '0';
    P14RI	: in std_logic := '0';
    P14RL	: in std_logic := '0';
    P14RR	: in std_logic := '0';
    P14RO1	: out std_logic := '0';
    P14RO2	: out std_logic := '0';
    P14RO3	: out std_logic := '0';
    P14RO4	: out std_logic := '0';
    P14RO5	: out std_logic := '0';

    P15CI1	: in std_logic := '0';
    P15CL	: in std_logic := '0';
    P15CR	: in std_logic := '0';
    P15CO	: out std_logic := '0';
    P15CTI	: in std_logic := '0';
    P15CTO	: out std_logic := '0';
    P15EI1	: in std_logic := '0';
    P15EI2	: in std_logic := '0';
    P15EI3	: in std_logic := '0';
    P15EI4	: in std_logic := '0';
    P15EI5	: in std_logic := '0';
    P15EL	: in std_logic := '0';
    P15ER	: in std_logic := '0';
    P15EO	: out std_logic := '0';
    P15RI	: in std_logic := '0';
    P15RL	: in std_logic := '0';
    P15RR	: in std_logic := '0';
    P15RO1	: out std_logic := '0';
    P15RO2	: out std_logic := '0';
    P15RO3	: out std_logic := '0';
    P15RO4	: out std_logic := '0';
    P15RO5	: out std_logic := '0';

    P16CI1	: in std_logic := '0';
    P16CL	: in std_logic := '0';
    P16CR	: in std_logic := '0';
    P16CO	: out std_logic := '0';
    P16CTI	: in std_logic := '0';
    P16CTO	: out std_logic := '0';
    P16EI1	: in std_logic := '0';
    P16EI2	: in std_logic := '0';
    P16EI3	: in std_logic := '0';
    P16EI4	: in std_logic := '0';
    P16EI5	: in std_logic := '0';
    P16EL	: in std_logic := '0';
    P16ER	: in std_logic := '0';
    P16EO	: out std_logic := '0';
    P16RI	: in std_logic := '0';
    P16RL	: in std_logic := '0';
    P16RR	: in std_logic := '0';
    P16RO1	: out std_logic := '0';
    P16RO2	: out std_logic := '0';
    P16RO3	: out std_logic := '0';
    P16RO4	: out std_logic := '0';
    P16RO5	: out std_logic := '0';

    P17CI1	: in std_logic := '0';
    P17CL	: in std_logic := '0';
    P17CR	: in std_logic := '0';
    P17CO	: out std_logic := '0';
    P17CTI	: in std_logic := '0';
    P17CTO	: out std_logic := '0';
    P17EI1	: in std_logic := '0';
    P17EI2	: in std_logic := '0';
    P17EI3	: in std_logic := '0';
    P17EI4	: in std_logic := '0';
    P17EI5	: in std_logic := '0';
    P17EL	: in std_logic := '0';
    P17ER	: in std_logic := '0';
    P17EO	: out std_logic := '0';
    P17RI	: in std_logic := '0';
    P17RL	: in std_logic := '0';
    P17RR	: in std_logic := '0';
    P17RO1	: out std_logic := '0';
    P17RO2	: out std_logic := '0';
    P17RO3	: out std_logic := '0';
    P17RO4	: out std_logic := '0';
    P17RO5	: out std_logic := '0';

    P18CI1	: in std_logic := '0';
    P18CL	: in std_logic := '0';
    P18CR	: in std_logic := '0';
    P18CO	: out std_logic := '0';
    P18CTI	: in std_logic := '0';
    P18CTO	: out std_logic := '0';
    P18EI1	: in std_logic := '0';
    P18EI2	: in std_logic := '0';
    P18EI3	: in std_logic := '0';
    P18EI4	: in std_logic := '0';
    P18EI5	: in std_logic := '0';
    P18EL	: in std_logic := '0';
    P18ER	: in std_logic := '0';
    P18EO	: out std_logic := '0';
    P18RI	: in std_logic := '0';
    P18RL	: in std_logic := '0';
    P18RR	: in std_logic := '0';
    P18RO1	: out std_logic := '0';
    P18RO2	: out std_logic := '0';
    P18RO3	: out std_logic := '0';
    P18RO4	: out std_logic := '0';
    P18RO5	: out std_logic := '0';

    P19CI1	: in std_logic := '0';
    P19CL	: in std_logic := '0';
    P19CR	: in std_logic := '0';
    P19CO	: out std_logic := '0';
    P19CTI	: in std_logic := '0';
    P19CTO	: out std_logic := '0';
    P19EI1	: in std_logic := '0';
    P19EI2	: in std_logic := '0';
    P19EI3	: in std_logic := '0';
    P19EI4	: in std_logic := '0';
    P19EI5	: in std_logic := '0';
    P19EL	: in std_logic := '0';
    P19ER	: in std_logic := '0';
    P19EO	: out std_logic := '0';
    P19RI	: in std_logic := '0';
    P19RL	: in std_logic := '0';
    P19RR	: in std_logic := '0';
    P19RO1	: out std_logic := '0';
    P19RO2	: out std_logic := '0';
    P19RO3	: out std_logic := '0';
    P19RO4	: out std_logic := '0';
    P19RO5	: out std_logic := '0';

    P20CI1	: in std_logic := '0';
    P20CL	: in std_logic := '0';
    P20CR	: in std_logic := '0';
    P20CO	: out std_logic := '0';
    P20CTI	: in std_logic := '0';
    P20CTO	: out std_logic := '0';
    P20EI1	: in std_logic := '0';
    P20EI2	: in std_logic := '0';
    P20EI3	: in std_logic := '0';
    P20EI4	: in std_logic := '0';
    P20EI5	: in std_logic := '0';
    P20EL	: in std_logic := '0';
    P20ER	: in std_logic := '0';
    P20EO	: out std_logic := '0';
    P20RI	: in std_logic := '0';
    P20RL	: in std_logic := '0';
    P20RR	: in std_logic := '0';
    P20RO1	: out std_logic := '0';
    P20RO2	: out std_logic := '0';
    P20RO3	: out std_logic := '0';
    P20RO4	: out std_logic := '0';
    P20RO5	: out std_logic := '0';

    P21CI1	: in std_logic := '0';
    P21CL	: in std_logic := '0';
    P21CR	: in std_logic := '0';
    P21CO	: out std_logic := '0';
    P21CTI	: in std_logic := '0';
    P21CTO	: out std_logic := '0';
    P21EI1	: in std_logic := '0';
    P21EI2	: in std_logic := '0';
    P21EI3	: in std_logic := '0';
    P21EI4	: in std_logic := '0';
    P21EI5	: in std_logic := '0';
    P21EL	: in std_logic := '0';
    P21ER	: in std_logic := '0';
    P21EO	: out std_logic := '0';
    P21RI	: in std_logic := '0';
    P21RL	: in std_logic := '0';
    P21RR	: in std_logic := '0';
    P21RO1	: out std_logic := '0';
    P21RO2	: out std_logic := '0';
    P21RO3	: out std_logic := '0';
    P21RO4	: out std_logic := '0';
    P21RO5	: out std_logic := '0';

    P22CI1	: in std_logic := '0';
    P22CL	: in std_logic := '0';
    P22CR	: in std_logic := '0';
    P22CO	: out std_logic := '0';
    P22CTI	: in std_logic := '0';
    P22CTO	: out std_logic := '0';
    P22EI1	: in std_logic := '0';
    P22EI2	: in std_logic := '0';
    P22EI3	: in std_logic := '0';
    P22EI4	: in std_logic := '0';
    P22EI5	: in std_logic := '0';
    P22EL	: in std_logic := '0';
    P22ER	: in std_logic := '0';
    P22EO	: out std_logic := '0';
    P22RI	: in std_logic := '0';
    P22RL	: in std_logic := '0';
    P22RR	: in std_logic := '0';
    P22RO1	: out std_logic := '0';
    P22RO2	: out std_logic := '0';
    P22RO3	: out std_logic := '0';
    P22RO4	: out std_logic := '0';
    P22RO5	: out std_logic := '0';

    P23CI1	: in std_logic := '0';
    P23CL	: in std_logic := '0';
    P23CR	: in std_logic := '0';
    P23CO	: out std_logic := '0';
    P23CTI	: in std_logic := '0';
    P23CTO	: out std_logic := '0';
    P23EI1	: in std_logic := '0';
    P23EI2	: in std_logic := '0';
    P23EI3	: in std_logic := '0';
    P23EI4	: in std_logic := '0';
    P23EI5	: in std_logic := '0';
    P23EL	: in std_logic := '0';
    P23ER	: in std_logic := '0';
    P23EO	: out std_logic := '0';
    P23RI	: in std_logic := '0';
    P23RL	: in std_logic := '0';
    P23RR	: in std_logic := '0';
    P23RO1	: out std_logic := '0';
    P23RO2	: out std_logic := '0';
    P23RO3	: out std_logic := '0';
    P23RO4	: out std_logic := '0';
    P23RO5	: out std_logic := '0';

    P24CI1	: in std_logic := '0';
    P24CL	: in std_logic := '0';
    P24CR	: in std_logic := '0';
    P24CO	: out std_logic := '0';
    P24CTI	: in std_logic := '0';
    P24CTO	: out std_logic := '0';
    P24EI1	: in std_logic := '0';
    P24EI2	: in std_logic := '0';
    P24EI3	: in std_logic := '0';
    P24EI4	: in std_logic := '0';
    P24EI5	: in std_logic := '0';
    P24EL	: in std_logic := '0';
    P24ER	: in std_logic := '0';
    P24EO	: out std_logic := '0';
    P24RI	: in std_logic := '0';
    P24RL	: in std_logic := '0';
    P24RR	: in std_logic := '0';
    P24RO1	: out std_logic := '0';
    P24RO2	: out std_logic := '0';
    P24RO3	: out std_logic := '0';
    P24RO4	: out std_logic := '0';
    P24RO5	: out std_logic := '0';

    P25CI1	: in std_logic := '0';
    P25CL	: in std_logic := '0';
    P25CR	: in std_logic := '0';
    P25CO	: out std_logic := '0';
    P25CTI	: in std_logic := '0';
    P25CTO	: out std_logic := '0';
    P25EI1	: in std_logic := '0';
    P25EI2	: in std_logic := '0';
    P25EI3	: in std_logic := '0';
    P25EI4	: in std_logic := '0';
    P25EI5	: in std_logic := '0';
    P25EL	: in std_logic := '0';
    P25ER	: in std_logic := '0';
    P25EO	: out std_logic := '0';
    P25RI	: in std_logic := '0';
    P25RL	: in std_logic := '0';
    P25RR	: in std_logic := '0';
    P25RO1	: out std_logic := '0';
    P25RO2	: out std_logic := '0';
    P25RO3	: out std_logic := '0';
    P25RO4	: out std_logic := '0';
    P25RO5	: out std_logic := '0';

    P26CI1	: in std_logic := '0';
    P26CL	: in std_logic := '0';
    P26CR	: in std_logic := '0';
    P26CO	: out std_logic := '0';
    P26CTI	: in std_logic := '0';
    P26CTO	: out std_logic := '0';
    P26EI1	: in std_logic := '0';
    P26EI2	: in std_logic := '0';
    P26EI3	: in std_logic := '0';
    P26EI4	: in std_logic := '0';
    P26EI5	: in std_logic := '0';
    P26EL	: in std_logic := '0';
    P26ER	: in std_logic := '0';
    P26EO	: out std_logic := '0';
    P26RI	: in std_logic := '0';
    P26RL	: in std_logic := '0';
    P26RR	: in std_logic := '0';
    P26RO1	: out std_logic := '0';
    P26RO2	: out std_logic := '0';
    P26RO3	: out std_logic := '0';
    P26RO4	: out std_logic := '0';
    P26RO5	: out std_logic := '0';

    P27CI1	: in std_logic := '0';
    P27CL	: in std_logic := '0';
    P27CR	: in std_logic := '0';
    P27CO	: out std_logic := '0';
    P27CTI	: in std_logic := '0';
    P27CTO	: out std_logic := '0';
    P27EI1	: in std_logic := '0';
    P27EI2	: in std_logic := '0';
    P27EI3	: in std_logic := '0';
    P27EI4	: in std_logic := '0';
    P27EI5	: in std_logic := '0';
    P27EL	: in std_logic := '0';
    P27ER	: in std_logic := '0';
    P27EO	: out std_logic := '0';
    P27RI	: in std_logic := '0';
    P27RL	: in std_logic := '0';
    P27RR	: in std_logic := '0';
    P27RO1	: out std_logic := '0';
    P27RO2	: out std_logic := '0';
    P27RO3	: out std_logic := '0';
    P27RO4	: out std_logic := '0';
    P27RO5	: out std_logic := '0';

    P28CI1	: in std_logic := '0';
    P28CL	: in std_logic := '0';
    P28CR	: in std_logic := '0';
    P28CO	: out std_logic := '0';
    P28CTI	: in std_logic := '0';
    P28CTO	: out std_logic := '0';
    P28EI1	: in std_logic := '0';
    P28EI2	: in std_logic := '0';
    P28EI3	: in std_logic := '0';
    P28EI4	: in std_logic := '0';
    P28EI5	: in std_logic := '0';
    P28EL	: in std_logic := '0';
    P28ER	: in std_logic := '0';
    P28EO	: out std_logic := '0';
    P28RI	: in std_logic := '0';
    P28RL	: in std_logic := '0';
    P28RR	: in std_logic := '0';
    P28RO1	: out std_logic := '0';
    P28RO2	: out std_logic := '0';
    P28RO3	: out std_logic := '0';
    P28RO4	: out std_logic := '0';
    P28RO5	: out std_logic := '0';

    P29CI1	: in std_logic := '0';
    P29CI2	: in std_logic := '0';
    P29CI3	: in std_logic := '0';
    P29CI4	: in std_logic := '0';
    P29CI5	: in std_logic := '0';
    P29CL	: in std_logic := '0';
    P29CR	: in std_logic := '0';
    P29CO	: out std_logic := '0';
    P29CTI	: in std_logic := '0';
    P29CTO	: out std_logic := '0';
    P29EI1	: in std_logic := '0';
    P29EI2	: in std_logic := '0';
    P29EI3	: in std_logic := '0';
    P29EI4	: in std_logic := '0';
    P29EI5	: in std_logic := '0';
    P29EL	: in std_logic := '0';
    P29ER	: in std_logic := '0';
    P29EO	: out std_logic := '0';
    P29RI	: in std_logic := '0';
    P29RL	: in std_logic := '0';
    P29RR	: in std_logic := '0';
    P29RO1	: out std_logic := '0';
    P29RO2	: out std_logic := '0';
    P29RO3	: out std_logic := '0';
    P29RO4	: out std_logic := '0';
    P29RO5	: out std_logic := '0';

    P30CI1	: in std_logic := '0';
    P30CL	: in std_logic := '0';
    P30CR	: in std_logic := '0';
    P30CO	: out std_logic := '0';
    P30CTI	: in std_logic := '0';
    P30CTO	: out std_logic := '0';
    P30EI1	: in std_logic := '0';
    P30EI2	: in std_logic := '0';
    P30EI3	: in std_logic := '0';
    P30EI4	: in std_logic := '0';
    P30EI5	: in std_logic := '0';
    P30EL	: in std_logic := '0';
    P30ER	: in std_logic := '0';
    P30EO	: out std_logic := '0';
    P30RI	: in std_logic := '0';
    P30RL	: in std_logic := '0';
    P30RR	: in std_logic := '0';
    P30RO1	: out std_logic := '0';
    P30RO2	: out std_logic := '0';
    P30RO3	: out std_logic := '0';
    P30RO4	: out std_logic := '0';
    P30RO5	: out std_logic := '0';

    P31CI1	: in std_logic := '0';
    P31CL	: in std_logic := '0';
    P31CR	: in std_logic := '0';
    P31CO	: out std_logic := '0';
    P31CTI	: in std_logic := '0';
    P31CTO	: out std_logic := '0';
    P31EI1	: in std_logic := '0';
    P31EI2	: in std_logic := '0';
    P31EI3	: in std_logic := '0';
    P31EI4	: in std_logic := '0';
    P31EI5	: in std_logic := '0';
    P31EL	: in std_logic := '0';
    P31ER	: in std_logic := '0';
    P31EO	: out std_logic := '0';
    P31RI	: in std_logic := '0';
    P31RL	: in std_logic := '0';
    P31RR	: in std_logic := '0';
    P31RO1	: out std_logic := '0';
    P31RO2	: out std_logic := '0';
    P31RO3	: out std_logic := '0';
    P31RO4	: out std_logic := '0';
    P31RO5	: out std_logic := '0';

    P32CI1	: in std_logic := '0';
    P32CL	: in std_logic := '0';
    P32CR	: in std_logic := '0';
    P32CO	: out std_logic := '0';
    P32CTI	: in std_logic := '0';
    P32CTO	: out std_logic := '0';
    P32EI1	: in std_logic := '0';
    P32EI2	: in std_logic := '0';
    P32EI3	: in std_logic := '0';
    P32EI4	: in std_logic := '0';
    P32EI5	: in std_logic := '0';
    P32EL	: in std_logic := '0';
    P32ER	: in std_logic := '0';
    P32EO	: out std_logic := '0';
    P32RI	: in std_logic := '0';
    P32RL	: in std_logic := '0';
    P32RR	: in std_logic := '0';
    P32RO1	: out std_logic := '0';
    P32RO2	: out std_logic := '0';
    P32RO3	: out std_logic := '0';
    P32RO4	: out std_logic := '0';
    P32RO5	: out std_logic := '0';

    P33CI1	: in std_logic := '0';
    P33CL	: in std_logic := '0';
    P33CR	: in std_logic := '0';
    P33CO	: out std_logic := '0';
    P33CTI	: in std_logic := '0';
    P33CTO	: out std_logic := '0';
    P33EI1	: in std_logic := '0';
    P33EI2	: in std_logic := '0';
    P33EI3	: in std_logic := '0';
    P33EI4	: in std_logic := '0';
    P33EI5	: in std_logic := '0';
    P33EL	: in std_logic := '0';
    P33ER	: in std_logic := '0';
    P33EO	: out std_logic := '0';
    P33RI	: in std_logic := '0';
    P33RL	: in std_logic := '0';
    P33RR	: in std_logic := '0';
    P33RO1	: out std_logic := '0';
    P33RO2	: out std_logic := '0';
    P33RO3	: out std_logic := '0';
    P33RO4	: out std_logic := '0';
    P33RO5	: out std_logic := '0';

    P34CI1	: in std_logic := '0';
    P34CL	: in std_logic := '0';
    P34CR	: in std_logic := '0';
    P34CO	: out std_logic := '0';
    P34CTI	: in std_logic := '0';
    P34CTO	: out std_logic := '0';
    P34EI1	: in std_logic := '0';
    P34EI2	: in std_logic := '0';
    P34EI3	: in std_logic := '0';
    P34EI4	: in std_logic := '0';
    P34EI5	: in std_logic := '0';
    P34EL	: in std_logic := '0';
    P34ER	: in std_logic := '0';
    P34EO	: out std_logic := '0';
    P34RI	: in std_logic := '0';
    P34RL	: in std_logic := '0';
    P34RR	: in std_logic := '0';
    P34RO1	: out std_logic := '0';
    P34RO2	: out std_logic := '0';
    P34RO3	: out std_logic := '0';
    P34RO4	: out std_logic := '0';
    P34RO5	: out std_logic := '0'
);
end component NX_IOM_L;

component NX_IOM_CONTROL_L is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port (
    RTCK1	: in std_logic := '0';
    RRCK1	: in std_logic := '0';
    WTCK1	: in std_logic := '0';
    WRCK1	: in std_logic := '0';
    RTCK2	: in std_logic := '0';
    RRCK2	: in std_logic := '0';
    WTCK2	: in std_logic := '0';
    WRCK2	: in std_logic := '0';
    CTCK	: in std_logic := '0';

    C1TW	: in std_logic := '0';
    C1TS	: in std_logic := '0';
    C1RW1	: in std_logic := '0';
    C1RW2	: in std_logic := '0';
    C1RW3	: in std_logic := '0';
    C1RNE	: in std_logic := '0';
    C1RS	: in std_logic := '0';
    C2TW	: in std_logic := '0';
    C2TS	: in std_logic := '0';
    C2RW1	: in std_logic := '0';
    C2RW2	: in std_logic := '0';
    C2RW3	: in std_logic := '0';
    C2RNE	: in std_logic := '0';
    C2RS	: in std_logic := '0';
    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';
    DC	: in std_logic := '0';
    CCK	: in std_logic := '0';
    DCK	: in std_logic := '0';
    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';
    DRA5	: in std_logic := '0';
    DRA6	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DOS	: in std_logic := '0';
    DOG	: in std_logic := '0';
    DIS	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DPAS	: in std_logic := '0';
    DPAG	: in std_logic := '0';
    DQSS	: in std_logic := '0';
    DQSG	: in std_logic := '0';
    DS1	: in std_logic := '0';
    DS2	: in std_logic := '0';
    CAD1	: in std_logic := '0';
    CAD2	: in std_logic := '0';
    CAD3	: in std_logic := '0';
    CAD4	: in std_logic := '0';
    CAD5	: in std_logic := '0';
    CAD6	: in std_logic := '0';
    CAP1	: in std_logic := '0';
    CAP2	: in std_logic := '0';
    CAP3	: in std_logic := '0';
    CAP4	: in std_logic := '0';
    CAN1	: in std_logic := '0';
    CAN2	: in std_logic := '0';
    CAN3	: in std_logic := '0';
    CAN4	: in std_logic := '0';
    CAT1	: in std_logic := '0';
    CAT2	: in std_logic := '0';
    CAT3	: in std_logic := '0';
    CAT4	: in std_logic := '0';
    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    C1RED	: out std_logic := '0';
    C2RED	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';
    CAL	: out std_logic := '0';

    LINK1	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK2	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK3	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK4	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK5	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK6	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK7	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK8	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK9	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK10	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK11	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK12	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK13	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK14	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK15	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK16	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK17	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK18	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK19	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK20	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK21	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK22	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK23	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK24	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK25	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK26	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK27	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK28	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK29	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK30	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK31	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK32	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK33	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK34	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_CONTROL_L;

component NX_IOM_DRIVER_M is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit_vector(1 downto 0) := "00";

    variant         : string := "";
    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1	: in std_logic := '0';
    EI2	: in std_logic := '0';
    EI3	: in std_logic := '0';
    EI4	: in std_logic := '0';
    EI5	: in std_logic := '0';
    EL	: in std_logic := '0';
    ER	: in std_logic := '0';
    CI1	: in std_logic := '0';
    CI2	: in std_logic := '0';
    CI3	: in std_logic := '0';
    CI4	: in std_logic := '0';
    CI5	: in std_logic := '0';
    CL	: in std_logic := '0';
    CR	: in std_logic := '0';
    CTI	: in std_logic := '0';
    RI	: in std_logic := '0';
    RL	: in std_logic := '0';
    RR	: in std_logic := '0';
    CO	: out std_logic := '0';
    EO	: out std_logic := '0';
    RO1	: out std_logic := '0';
    RO2	: out std_logic := '0';
    RO3	: out std_logic := '0';
    RO4	: out std_logic := '0';
    RO5	: out std_logic := '0';
    CTO	: out std_logic := '0';
    LINK	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_DRIVER_M;

component NX_IOM_SERDES_M is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    RTCK	: in std_logic := '0';
    WRCK	: in std_logic := '0';
    WTCK	: in std_logic := '0';
    RRCK	: in std_logic := '0';
    TRST	: in std_logic := '0';
    RRST	: in std_logic := '0';
    CTCK	: in std_logic := '0';
    DCK	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DS	: in std_logic_vector(1 downto 0) := (others => '0');
    DRA	: in std_logic_vector(5 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');
    FZ	: in std_logic := '0';
    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0');
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    LINKN	: inout std_logic_vector(IOM_LINK_SIZE-1 downto 0) := (others => '0');
    LINKP	: inout std_logic_vector(IOM_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_IOM_SERDES_M;

component NX_IOM_DRIVER is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit_vector(1 downto 0) := "00";

    variant         : string := "";
    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1	: in std_logic := '0';
    EI2	: in std_logic := '0';
    EI3	: in std_logic := '0';
    EI4	: in std_logic := '0';
    EI5	: in std_logic := '0';
    EL	: in std_logic := '0';
    ER	: in std_logic := '0';
    CI1	: in std_logic := '0';
    CI2	: in std_logic := '0';
    CI3	: in std_logic := '0';
    CI4	: in std_logic := '0';
    CI5	: in std_logic := '0';
    CL	: in std_logic := '0';
    CR	: in std_logic := '0';
    CTI	: in std_logic := '0';
    RI	: in std_logic := '0';
    RL	: in std_logic := '0';
    RR	: in std_logic := '0';
    CO	: out std_logic := '0';
    EO	: out std_logic := '0';
    RO1	: out std_logic := '0';
    RO2	: out std_logic := '0';
    RO3	: out std_logic := '0';
    RO4	: out std_logic := '0';
    RO5	: out std_logic := '0';
    CTO	: out std_logic := '0';
    LINK	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_DRIVER;

component NX_IOM_CONTROL is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port (
    RTCK1	: in std_logic := '0';
    RRCK1	: in std_logic := '0';
    WTCK1	: in std_logic := '0';
    WRCK1	: in std_logic := '0';
    RTCK2	: in std_logic := '0';
    RRCK2	: in std_logic := '0';
    WTCK2	: in std_logic := '0';
    WRCK2	: in std_logic := '0';
    CTCK	: in std_logic := '0';

    C1TW	: in std_logic := '0';
    C1TS	: in std_logic := '0';
    C1RW1	: in std_logic := '0';
    C1RW2	: in std_logic := '0';
    C1RW3	: in std_logic := '0';
    C1RNE	: in std_logic := '0';
    C1RS	: in std_logic := '0';
    C2TW	: in std_logic := '0';
    C2TS	: in std_logic := '0';
    C2RW1	: in std_logic := '0';
    C2RW2	: in std_logic := '0';
    C2RW3	: in std_logic := '0';
    C2RNE	: in std_logic := '0';
    C2RS	: in std_logic := '0';
    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';
    DC	: in std_logic := '0';
    CCK	: in std_logic := '0';
    DCK	: in std_logic := '0';
    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';
    DRA5	: in std_logic := '0';
    DRA6	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DOS	: in std_logic := '0';
    DOG	: in std_logic := '0';
    DIS	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DPAS	: in std_logic := '0';
    DPAG	: in std_logic := '0';
    DQSS	: in std_logic := '0';
    DQSG	: in std_logic := '0';
    DS1	: in std_logic := '0';
    DS2	: in std_logic := '0';
    CAD1	: in std_logic := '0';
    CAD2	: in std_logic := '0';
    CAD3	: in std_logic := '0';
    CAD4	: in std_logic := '0';
    CAD5	: in std_logic := '0';
    CAD6	: in std_logic := '0';
    CAP1	: in std_logic := '0';
    CAP2	: in std_logic := '0';
    CAP3	: in std_logic := '0';
    CAP4	: in std_logic := '0';
    CAN1	: in std_logic := '0';
    CAN2	: in std_logic := '0';
    CAN3	: in std_logic := '0';
    CAN4	: in std_logic := '0';
    CAT1	: in std_logic := '0';
    CAT2	: in std_logic := '0';
    CAT3	: in std_logic := '0';
    CAT4	: in std_logic := '0';
    SPI1	: in std_logic := '0';
    SPI2	: in std_logic := '0';
    SPI3	: in std_logic := '0';
    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    C1RED	: out std_logic := '0';
    C2RED	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';
    CAL	: out std_logic := '0';

    LINK1	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK2	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK3	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK4	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK5	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK6	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK7	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK8	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK9	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK10	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK11	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK12	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK13	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK14	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK15	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK16	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK17	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK18	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK19	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK20	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK21	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK22	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK23	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK24	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK25	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK26	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK27	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK28	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK29	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK30	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK31	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK32	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK33	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK34	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_CONTROL;

component NX_IOM_SERDES is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    RTCK	: in std_logic := '0';
    WRCK	: in std_logic := '0';
    WTCK	: in std_logic := '0';
    RRCK	: in std_logic := '0';
    TRST	: in std_logic := '0';
    RRST	: in std_logic := '0';
    CTCK	: in std_logic := '0';
    DCK	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DS	: in std_logic_vector(1 downto 0) := (others => '0');
    DRA	: in std_logic_vector(5 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');
    FZ	: in std_logic := '0';
    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0');
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    LINKN	: inout std_logic_vector(IOM_LINK_SIZE-1 downto 0) := (others => '0');
    LINKP	: inout std_logic_vector(IOM_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_IOM_SERDES;

component NX_IOM is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk1 : bit := '0';
--  latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk2 : bit := '0';
--  latency2     : bit := '0';
--  sel_clk_out2 : bit_vector(1 downto 0) := "00";
--  sel_clk_out3 : bit_vector(1 downto 0) := "00";
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_io_cal  : bit := '0';
    pads_dict    : string := "";
    pads_path    : string := ""
);
port (
    RTCK1	: in std_logic := '0';
    RRCK1	: in std_logic := '0';
    WTCK1	: in std_logic := '0';
    WRCK1	: in std_logic := '0';
    RTCK2	: in std_logic := '0';
    RRCK2	: in std_logic := '0';
    WTCK2	: in std_logic := '0';
    WRCK2	: in std_logic := '0';
    CTCK	: in std_logic := '0';
    CCK	: in std_logic := '0';
    DCK	: in std_logic := '0';

    C1TW	: in std_logic := '0';
    C1TS	: in std_logic := '0';
    C1RW1	: in std_logic := '0';
    C1RW2	: in std_logic := '0';
    C1RW3	: in std_logic := '0';
    C1RNE	: in std_logic := '0';
    C1RS	: in std_logic := '0';
    C2TW	: in std_logic := '0';
    C2TS	: in std_logic := '0';
    C2RW1	: in std_logic := '0';
    C2RW2	: in std_logic := '0';
    C2RW3	: in std_logic := '0';
    C2RNE	: in std_logic := '0';
    C2RS	: in std_logic := '0';
    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FZ	: in std_logic := '0';
    DC	: in std_logic := '0';
    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';
    DRA5	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DOS	: in std_logic := '0';
    DOG	: in std_logic := '0';
    DIS	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DPAS	: in std_logic := '0';
    DPAG	: in std_logic := '0';
    DQSS	: in std_logic := '0';
    DQSG	: in std_logic := '0';
    DS1	: in std_logic := '0';
    DS2	: in std_logic := '0';
    CAD1	: in std_logic := '0';
    CAD2	: in std_logic := '0';
    CAD3	: in std_logic := '0';
    CAD4	: in std_logic := '0';
    CAD5	: in std_logic := '0';
    CAD6	: in std_logic := '0';
    CAP1	: in std_logic := '0';
    CAP2	: in std_logic := '0';
    CAP3	: in std_logic := '0';
    CAP4	: in std_logic := '0';
    CAN1	: in std_logic := '0';
    CAN2	: in std_logic := '0';
    CAN3	: in std_logic := '0';
    CAN4	: in std_logic := '0';
    CAT1	: in std_logic := '0';
    CAT2	: in std_logic := '0';
    CAT3	: in std_logic := '0';
    CAT4	: in std_logic := '0';
    SPI1	: in std_logic := '0';
    SPI2	: in std_logic := '0';
    SPI3	: in std_logic := '0';

    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';

    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    C1RED	: out std_logic := '0';
    C2RED	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';
    CAL	: out std_logic := '0';

    P1CI1	: in std_logic := '0';
    P1CL	: in std_logic := '0';
    P1CR	: in std_logic := '0';
    P1CO	: out std_logic := '0';
    P1CTI	: in std_logic := '0';
    P1CTO	: out std_logic := '0';
    P1EI1	: in std_logic := '0';
    P1EI2	: in std_logic := '0';
    P1EI3	: in std_logic := '0';
    P1EI4	: in std_logic := '0';
    P1EI5	: in std_logic := '0';
    P1EL	: in std_logic := '0';
    P1ER	: in std_logic := '0';
    P1EO	: out std_logic := '0';
    P1RI	: in std_logic := '0';
    P1RL	: in std_logic := '0';
    P1RR	: in std_logic := '0';
    P1RO1	: out std_logic := '0';
    P1RO2	: out std_logic := '0';
    P1RO3	: out std_logic := '0';
    P1RO4	: out std_logic := '0';
    P1RO5	: out std_logic := '0';

    P2CI1	: in std_logic := '0';
    P2CL	: in std_logic := '0';
    P2CR	: in std_logic := '0';
    P2CO	: out std_logic := '0';
    P2CTI	: in std_logic := '0';
    P2CTO	: out std_logic := '0';
    P2EI1	: in std_logic := '0';
    P2EI2	: in std_logic := '0';
    P2EI3	: in std_logic := '0';
    P2EI4	: in std_logic := '0';
    P2EI5	: in std_logic := '0';
    P2EL	: in std_logic := '0';
    P2ER	: in std_logic := '0';
    P2EO	: out std_logic := '0';
    P2RI	: in std_logic := '0';
    P2RL	: in std_logic := '0';
    P2RR	: in std_logic := '0';
    P2RO1	: out std_logic := '0';
    P2RO2	: out std_logic := '0';
    P2RO3	: out std_logic := '0';
    P2RO4	: out std_logic := '0';
    P2RO5	: out std_logic := '0';

    P3CI1	: in std_logic := '0';
    P3CL	: in std_logic := '0';
    P3CR	: in std_logic := '0';
    P3CO	: out std_logic := '0';
    P3CTI	: in std_logic := '0';
    P3CTO	: out std_logic := '0';
    P3EI1	: in std_logic := '0';
    P3EI2	: in std_logic := '0';
    P3EI3	: in std_logic := '0';
    P3EI4	: in std_logic := '0';
    P3EI5	: in std_logic := '0';
    P3EL	: in std_logic := '0';
    P3ER	: in std_logic := '0';
    P3EO	: out std_logic := '0';
    P3RI	: in std_logic := '0';
    P3RL	: in std_logic := '0';
    P3RR	: in std_logic := '0';
    P3RO1	: out std_logic := '0';
    P3RO2	: out std_logic := '0';
    P3RO3	: out std_logic := '0';
    P3RO4	: out std_logic := '0';
    P3RO5	: out std_logic := '0';

    P4CI1	: in std_logic := '0';
    P4CL	: in std_logic := '0';
    P4CR	: in std_logic := '0';
    P4CO	: out std_logic := '0';
    P4CTI	: in std_logic := '0';
    P4CTO	: out std_logic := '0';
    P4EI1	: in std_logic := '0';
    P4EI2	: in std_logic := '0';
    P4EI3	: in std_logic := '0';
    P4EI4	: in std_logic := '0';
    P4EI5	: in std_logic := '0';
    P4EL	: in std_logic := '0';
    P4ER	: in std_logic := '0';
    P4EO	: out std_logic := '0';
    P4RI	: in std_logic := '0';
    P4RL	: in std_logic := '0';
    P4RR	: in std_logic := '0';
    P4RO1	: out std_logic := '0';
    P4RO2	: out std_logic := '0';
    P4RO3	: out std_logic := '0';
    P4RO4	: out std_logic := '0';
    P4RO5	: out std_logic := '0';

    P5CI1	: in std_logic := '0';
    P5CI2	: in std_logic := '0';
    P5CI3	: in std_logic := '0';
    P5CI4	: in std_logic := '0';
    P5CI5	: in std_logic := '0';
    P5CL	: in std_logic := '0';
    P5CR	: in std_logic := '0';
    P5CO	: out std_logic := '0';
    P5CTI	: in std_logic := '0';
    P5CTO	: out std_logic := '0';
    P5EI1	: in std_logic := '0';
    P5EI2	: in std_logic := '0';
    P5EI3	: in std_logic := '0';
    P5EI4	: in std_logic := '0';
    P5EI5	: in std_logic := '0';
    P5EL	: in std_logic := '0';
    P5ER	: in std_logic := '0';
    P5EO	: out std_logic := '0';
    P5RI	: in std_logic := '0';
    P5RL	: in std_logic := '0';
    P5RR	: in std_logic := '0';
    P5RO1	: out std_logic := '0';
    P5RO2	: out std_logic := '0';
    P5RO3	: out std_logic := '0';
    P5RO4	: out std_logic := '0';
    P5RO5	: out std_logic := '0';

    P6CI1	: in std_logic := '0';
    P6CL	: in std_logic := '0';
    P6CR	: in std_logic := '0';
    P6CO	: out std_logic := '0';
    P6CTI	: in std_logic := '0';
    P6CTO	: out std_logic := '0';
    P6EI1	: in std_logic := '0';
    P6EI2	: in std_logic := '0';
    P6EI3	: in std_logic := '0';
    P6EI4	: in std_logic := '0';
    P6EI5	: in std_logic := '0';
    P6EL	: in std_logic := '0';
    P6ER	: in std_logic := '0';
    P6EO	: out std_logic := '0';
    P6RI	: in std_logic := '0';
    P6RL	: in std_logic := '0';
    P6RR	: in std_logic := '0';
    P6RO1	: out std_logic := '0';
    P6RO2	: out std_logic := '0';
    P6RO3	: out std_logic := '0';
    P6RO4	: out std_logic := '0';
    P6RO5	: out std_logic := '0';

    P7CI1	: in std_logic := '0';
    P7CL	: in std_logic := '0';
    P7CR	: in std_logic := '0';
    P7CO	: out std_logic := '0';
    P7CTI	: in std_logic := '0';
    P7CTO	: out std_logic := '0';
    P7EI1	: in std_logic := '0';
    P7EI2	: in std_logic := '0';
    P7EI3	: in std_logic := '0';
    P7EI4	: in std_logic := '0';
    P7EI5	: in std_logic := '0';
    P7EL	: in std_logic := '0';
    P7ER	: in std_logic := '0';
    P7EO	: out std_logic := '0';
    P7RI	: in std_logic := '0';
    P7RL	: in std_logic := '0';
    P7RR	: in std_logic := '0';
    P7RO1	: out std_logic := '0';
    P7RO2	: out std_logic := '0';
    P7RO3	: out std_logic := '0';
    P7RO4	: out std_logic := '0';
    P7RO5	: out std_logic := '0';

    P8CI1	: in std_logic := '0';
    P8CL	: in std_logic := '0';
    P8CR	: in std_logic := '0';
    P8CO	: out std_logic := '0';
    P8CTI	: in std_logic := '0';
    P8CTO	: out std_logic := '0';
    P8EI1	: in std_logic := '0';
    P8EI2	: in std_logic := '0';
    P8EI3	: in std_logic := '0';
    P8EI4	: in std_logic := '0';
    P8EI5	: in std_logic := '0';
    P8EL	: in std_logic := '0';
    P8ER	: in std_logic := '0';
    P8EO	: out std_logic := '0';
    P8RI	: in std_logic := '0';
    P8RL	: in std_logic := '0';
    P8RR	: in std_logic := '0';
    P8RO1	: out std_logic := '0';
    P8RO2	: out std_logic := '0';
    P8RO3	: out std_logic := '0';
    P8RO4	: out std_logic := '0';
    P8RO5	: out std_logic := '0';

    P9CI1	: in std_logic := '0';
    P9CL	: in std_logic := '0';
    P9CR	: in std_logic := '0';
    P9CO	: out std_logic := '0';
    P9CTI	: in std_logic := '0';
    P9CTO	: out std_logic := '0';
    P9EI1	: in std_logic := '0';
    P9EI2	: in std_logic := '0';
    P9EI3	: in std_logic := '0';
    P9EI4	: in std_logic := '0';
    P9EI5	: in std_logic := '0';
    P9EL	: in std_logic := '0';
    P9ER	: in std_logic := '0';
    P9EO	: out std_logic := '0';
    P9RI	: in std_logic := '0';
    P9RL	: in std_logic := '0';
    P9RR	: in std_logic := '0';
    P9RO1	: out std_logic := '0';
    P9RO2	: out std_logic := '0';
    P9RO3	: out std_logic := '0';
    P9RO4	: out std_logic := '0';
    P9RO5	: out std_logic := '0';

    P10CI1	: in std_logic := '0';
    P10CL	: in std_logic := '0';
    P10CR	: in std_logic := '0';
    P10CO	: out std_logic := '0';
    P10CTI	: in std_logic := '0';
    P10CTO	: out std_logic := '0';
    P10EI1	: in std_logic := '0';
    P10EI2	: in std_logic := '0';
    P10EI3	: in std_logic := '0';
    P10EI4	: in std_logic := '0';
    P10EI5	: in std_logic := '0';
    P10EL	: in std_logic := '0';
    P10ER	: in std_logic := '0';
    P10EO	: out std_logic := '0';
    P10RI	: in std_logic := '0';
    P10RL	: in std_logic := '0';
    P10RR	: in std_logic := '0';
    P10RO1	: out std_logic := '0';
    P10RO2	: out std_logic := '0';
    P10RO3	: out std_logic := '0';
    P10RO4	: out std_logic := '0';
    P10RO5	: out std_logic := '0';

    P11CI1	: in std_logic := '0';
    P11CL	: in std_logic := '0';
    P11CR	: in std_logic := '0';
    P11CO	: out std_logic := '0';
    P11CTI	: in std_logic := '0';
    P11CTO	: out std_logic := '0';
    P11EI1	: in std_logic := '0';
    P11EI2	: in std_logic := '0';
    P11EI3	: in std_logic := '0';
    P11EI4	: in std_logic := '0';
    P11EI5	: in std_logic := '0';
    P11EL	: in std_logic := '0';
    P11ER	: in std_logic := '0';
    P11EO	: out std_logic := '0';
    P11RI	: in std_logic := '0';
    P11RL	: in std_logic := '0';
    P11RR	: in std_logic := '0';
    P11RO1	: out std_logic := '0';
    P11RO2	: out std_logic := '0';
    P11RO3	: out std_logic := '0';
    P11RO4	: out std_logic := '0';
    P11RO5	: out std_logic := '0';

    P12CI1	: in std_logic := '0';
    P12CL	: in std_logic := '0';
    P12CR	: in std_logic := '0';
    P12CO	: out std_logic := '0';
    P12CTI	: in std_logic := '0';
    P12CTO	: out std_logic := '0';
    P12EI1	: in std_logic := '0';
    P12EI2	: in std_logic := '0';
    P12EI3	: in std_logic := '0';
    P12EI4	: in std_logic := '0';
    P12EI5	: in std_logic := '0';
    P12EL	: in std_logic := '0';
    P12ER	: in std_logic := '0';
    P12EO	: out std_logic := '0';
    P12RI	: in std_logic := '0';
    P12RL	: in std_logic := '0';
    P12RR	: in std_logic := '0';
    P12RO1	: out std_logic := '0';
    P12RO2	: out std_logic := '0';
    P12RO3	: out std_logic := '0';
    P12RO4	: out std_logic := '0';
    P12RO5	: out std_logic := '0';

    P13CI1	: in std_logic := '0';
    P13CL	: in std_logic := '0';
    P13CR	: in std_logic := '0';
    P13CO	: out std_logic := '0';
    P13CTI	: in std_logic := '0';
    P13CTO	: out std_logic := '0';
    P13EI1	: in std_logic := '0';
    P13EI2	: in std_logic := '0';
    P13EI3	: in std_logic := '0';
    P13EI4	: in std_logic := '0';
    P13EI5	: in std_logic := '0';
    P13EL	: in std_logic := '0';
    P13ER	: in std_logic := '0';
    P13EO	: out std_logic := '0';
    P13RI	: in std_logic := '0';
    P13RL	: in std_logic := '0';
    P13RR	: in std_logic := '0';
    P13RO1	: out std_logic := '0';
    P13RO2	: out std_logic := '0';
    P13RO3	: out std_logic := '0';
    P13RO4	: out std_logic := '0';
    P13RO5	: out std_logic := '0';

    P14CI1	: in std_logic := '0';
    P14CL	: in std_logic := '0';
    P14CR	: in std_logic := '0';
    P14CO	: out std_logic := '0';
    P14CTI	: in std_logic := '0';
    P14CTO	: out std_logic := '0';
    P14EI1	: in std_logic := '0';
    P14EI2	: in std_logic := '0';
    P14EI3	: in std_logic := '0';
    P14EI4	: in std_logic := '0';
    P14EI5	: in std_logic := '0';
    P14EL	: in std_logic := '0';
    P14ER	: in std_logic := '0';
    P14EO	: out std_logic := '0';
    P14RI	: in std_logic := '0';
    P14RL	: in std_logic := '0';
    P14RR	: in std_logic := '0';
    P14RO1	: out std_logic := '0';
    P14RO2	: out std_logic := '0';
    P14RO3	: out std_logic := '0';
    P14RO4	: out std_logic := '0';
    P14RO5	: out std_logic := '0';

    P15CI1	: in std_logic := '0';
    P15CL	: in std_logic := '0';
    P15CR	: in std_logic := '0';
    P15CO	: out std_logic := '0';
    P15CTI	: in std_logic := '0';
    P15CTO	: out std_logic := '0';
    P15EI1	: in std_logic := '0';
    P15EI2	: in std_logic := '0';
    P15EI3	: in std_logic := '0';
    P15EI4	: in std_logic := '0';
    P15EI5	: in std_logic := '0';
    P15EL	: in std_logic := '0';
    P15ER	: in std_logic := '0';
    P15EO	: out std_logic := '0';
    P15RI	: in std_logic := '0';
    P15RL	: in std_logic := '0';
    P15RR	: in std_logic := '0';
    P15RO1	: out std_logic := '0';
    P15RO2	: out std_logic := '0';
    P15RO3	: out std_logic := '0';
    P15RO4	: out std_logic := '0';
    P15RO5	: out std_logic := '0';

    P16CI1	: in std_logic := '0';
    P16CL	: in std_logic := '0';
    P16CR	: in std_logic := '0';
    P16CO	: out std_logic := '0';
    P16CTI	: in std_logic := '0';
    P16CTO	: out std_logic := '0';
    P16EI1	: in std_logic := '0';
    P16EI2	: in std_logic := '0';
    P16EI3	: in std_logic := '0';
    P16EI4	: in std_logic := '0';
    P16EI5	: in std_logic := '0';
    P16EL	: in std_logic := '0';
    P16ER	: in std_logic := '0';
    P16EO	: out std_logic := '0';
    P16RI	: in std_logic := '0';
    P16RL	: in std_logic := '0';
    P16RR	: in std_logic := '0';
    P16RO1	: out std_logic := '0';
    P16RO2	: out std_logic := '0';
    P16RO3	: out std_logic := '0';
    P16RO4	: out std_logic := '0';
    P16RO5	: out std_logic := '0';

    P17CI1	: in std_logic := '0';
    P17CL	: in std_logic := '0';
    P17CR	: in std_logic := '0';
    P17CO	: out std_logic := '0';
    P17CTI	: in std_logic := '0';
    P17CTO	: out std_logic := '0';
    P17EI1	: in std_logic := '0';
    P17EI2	: in std_logic := '0';
    P17EI3	: in std_logic := '0';
    P17EI4	: in std_logic := '0';
    P17EI5	: in std_logic := '0';
    P17EL	: in std_logic := '0';
    P17ER	: in std_logic := '0';
    P17EO	: out std_logic := '0';
    P17RI	: in std_logic := '0';
    P17RL	: in std_logic := '0';
    P17RR	: in std_logic := '0';
    P17RO1	: out std_logic := '0';
    P17RO2	: out std_logic := '0';
    P17RO3	: out std_logic := '0';
    P17RO4	: out std_logic := '0';
    P17RO5	: out std_logic := '0';

    P18CI1	: in std_logic := '0';
    P18CL	: in std_logic := '0';
    P18CR	: in std_logic := '0';
    P18CO	: out std_logic := '0';
    P18CTI	: in std_logic := '0';
    P18CTO	: out std_logic := '0';
    P18EI1	: in std_logic := '0';
    P18EI2	: in std_logic := '0';
    P18EI3	: in std_logic := '0';
    P18EI4	: in std_logic := '0';
    P18EI5	: in std_logic := '0';
    P18EL	: in std_logic := '0';
    P18ER	: in std_logic := '0';
    P18EO	: out std_logic := '0';
    P18RI	: in std_logic := '0';
    P18RL	: in std_logic := '0';
    P18RR	: in std_logic := '0';
    P18RO1	: out std_logic := '0';
    P18RO2	: out std_logic := '0';
    P18RO3	: out std_logic := '0';
    P18RO4	: out std_logic := '0';
    P18RO5	: out std_logic := '0';

    P19CI1	: in std_logic := '0';
    P19CL	: in std_logic := '0';
    P19CR	: in std_logic := '0';
    P19CO	: out std_logic := '0';
    P19CTI	: in std_logic := '0';
    P19CTO	: out std_logic := '0';
    P19EI1	: in std_logic := '0';
    P19EI2	: in std_logic := '0';
    P19EI3	: in std_logic := '0';
    P19EI4	: in std_logic := '0';
    P19EI5	: in std_logic := '0';
    P19EL	: in std_logic := '0';
    P19ER	: in std_logic := '0';
    P19EO	: out std_logic := '0';
    P19RI	: in std_logic := '0';
    P19RL	: in std_logic := '0';
    P19RR	: in std_logic := '0';
    P19RO1	: out std_logic := '0';
    P19RO2	: out std_logic := '0';
    P19RO3	: out std_logic := '0';
    P19RO4	: out std_logic := '0';
    P19RO5	: out std_logic := '0';

    P20CI1	: in std_logic := '0';
    P20CL	: in std_logic := '0';
    P20CR	: in std_logic := '0';
    P20CO	: out std_logic := '0';
    P20CTI	: in std_logic := '0';
    P20CTO	: out std_logic := '0';
    P20EI1	: in std_logic := '0';
    P20EI2	: in std_logic := '0';
    P20EI3	: in std_logic := '0';
    P20EI4	: in std_logic := '0';
    P20EI5	: in std_logic := '0';
    P20EL	: in std_logic := '0';
    P20ER	: in std_logic := '0';
    P20EO	: out std_logic := '0';
    P20RI	: in std_logic := '0';
    P20RL	: in std_logic := '0';
    P20RR	: in std_logic := '0';
    P20RO1	: out std_logic := '0';
    P20RO2	: out std_logic := '0';
    P20RO3	: out std_logic := '0';
    P20RO4	: out std_logic := '0';
    P20RO5	: out std_logic := '0';

    P21CI1	: in std_logic := '0';
    P21CL	: in std_logic := '0';
    P21CR	: in std_logic := '0';
    P21CO	: out std_logic := '0';
    P21CTI	: in std_logic := '0';
    P21CTO	: out std_logic := '0';
    P21EI1	: in std_logic := '0';
    P21EI2	: in std_logic := '0';
    P21EI3	: in std_logic := '0';
    P21EI4	: in std_logic := '0';
    P21EI5	: in std_logic := '0';
    P21EL	: in std_logic := '0';
    P21ER	: in std_logic := '0';
    P21EO	: out std_logic := '0';
    P21RI	: in std_logic := '0';
    P21RL	: in std_logic := '0';
    P21RR	: in std_logic := '0';
    P21RO1	: out std_logic := '0';
    P21RO2	: out std_logic := '0';
    P21RO3	: out std_logic := '0';
    P21RO4	: out std_logic := '0';
    P21RO5	: out std_logic := '0';

    P22CI1	: in std_logic := '0';
    P22CL	: in std_logic := '0';
    P22CR	: in std_logic := '0';
    P22CO	: out std_logic := '0';
    P22CTI	: in std_logic := '0';
    P22CTO	: out std_logic := '0';
    P22EI1	: in std_logic := '0';
    P22EI2	: in std_logic := '0';
    P22EI3	: in std_logic := '0';
    P22EI4	: in std_logic := '0';
    P22EI5	: in std_logic := '0';
    P22EL	: in std_logic := '0';
    P22ER	: in std_logic := '0';
    P22EO	: out std_logic := '0';
    P22RI	: in std_logic := '0';
    P22RL	: in std_logic := '0';
    P22RR	: in std_logic := '0';
    P22RO1	: out std_logic := '0';
    P22RO2	: out std_logic := '0';
    P22RO3	: out std_logic := '0';
    P22RO4	: out std_logic := '0';
    P22RO5	: out std_logic := '0';

    P23CI1	: in std_logic := '0';
    P23CL	: in std_logic := '0';
    P23CR	: in std_logic := '0';
    P23CO	: out std_logic := '0';
    P23CTI	: in std_logic := '0';
    P23CTO	: out std_logic := '0';
    P23EI1	: in std_logic := '0';
    P23EI2	: in std_logic := '0';
    P23EI3	: in std_logic := '0';
    P23EI4	: in std_logic := '0';
    P23EI5	: in std_logic := '0';
    P23EL	: in std_logic := '0';
    P23ER	: in std_logic := '0';
    P23EO	: out std_logic := '0';
    P23RI	: in std_logic := '0';
    P23RL	: in std_logic := '0';
    P23RR	: in std_logic := '0';
    P23RO1	: out std_logic := '0';
    P23RO2	: out std_logic := '0';
    P23RO3	: out std_logic := '0';
    P23RO4	: out std_logic := '0';
    P23RO5	: out std_logic := '0';

    P24CI1	: in std_logic := '0';
    P24CL	: in std_logic := '0';
    P24CR	: in std_logic := '0';
    P24CO	: out std_logic := '0';
    P24CTI	: in std_logic := '0';
    P24CTO	: out std_logic := '0';
    P24EI1	: in std_logic := '0';
    P24EI2	: in std_logic := '0';
    P24EI3	: in std_logic := '0';
    P24EI4	: in std_logic := '0';
    P24EI5	: in std_logic := '0';
    P24EL	: in std_logic := '0';
    P24ER	: in std_logic := '0';
    P24EO	: out std_logic := '0';
    P24RI	: in std_logic := '0';
    P24RL	: in std_logic := '0';
    P24RR	: in std_logic := '0';
    P24RO1	: out std_logic := '0';
    P24RO2	: out std_logic := '0';
    P24RO3	: out std_logic := '0';
    P24RO4	: out std_logic := '0';
    P24RO5	: out std_logic := '0';

    P25CI1	: in std_logic := '0';
    P25CI2	: in std_logic := '0';
    P25CI3	: in std_logic := '0';
    P25CI4	: in std_logic := '0';
    P25CI5	: in std_logic := '0';
    P25CL	: in std_logic := '0';
    P25CR	: in std_logic := '0';
    P25CO	: out std_logic := '0';
    P25CTI	: in std_logic := '0';
    P25CTO	: out std_logic := '0';
    P25EI1	: in std_logic := '0';
    P25EI2	: in std_logic := '0';
    P25EI3	: in std_logic := '0';
    P25EI4	: in std_logic := '0';
    P25EI5	: in std_logic := '0';
    P25EL	: in std_logic := '0';
    P25ER	: in std_logic := '0';
    P25EO	: out std_logic := '0';
    P25RI	: in std_logic := '0';
    P25RL	: in std_logic := '0';
    P25RR	: in std_logic := '0';
    P25RO1	: out std_logic := '0';
    P25RO2	: out std_logic := '0';
    P25RO3	: out std_logic := '0';
    P25RO4	: out std_logic := '0';
    P25RO5	: out std_logic := '0';

    P26CI1	: in std_logic := '0';
    P26CL	: in std_logic := '0';
    P26CR	: in std_logic := '0';
    P26CO	: out std_logic := '0';
    P26CTI	: in std_logic := '0';
    P26CTO	: out std_logic := '0';
    P26EI1	: in std_logic := '0';
    P26EI2	: in std_logic := '0';
    P26EI3	: in std_logic := '0';
    P26EI4	: in std_logic := '0';
    P26EI5	: in std_logic := '0';
    P26EL	: in std_logic := '0';
    P26ER	: in std_logic := '0';
    P26EO	: out std_logic := '0';
    P26RI	: in std_logic := '0';
    P26RL	: in std_logic := '0';
    P26RR	: in std_logic := '0';
    P26RO1	: out std_logic := '0';
    P26RO2	: out std_logic := '0';
    P26RO3	: out std_logic := '0';
    P26RO4	: out std_logic := '0';
    P26RO5	: out std_logic := '0';

    P27CI1	: in std_logic := '0';
    P27CL	: in std_logic := '0';
    P27CR	: in std_logic := '0';
    P27CO	: out std_logic := '0';
    P27CTI	: in std_logic := '0';
    P27CTO	: out std_logic := '0';
    P27EI1	: in std_logic := '0';
    P27EI2	: in std_logic := '0';
    P27EI3	: in std_logic := '0';
    P27EI4	: in std_logic := '0';
    P27EI5	: in std_logic := '0';
    P27EL	: in std_logic := '0';
    P27ER	: in std_logic := '0';
    P27EO	: out std_logic := '0';
    P27RI	: in std_logic := '0';
    P27RL	: in std_logic := '0';
    P27RR	: in std_logic := '0';
    P27RO1	: out std_logic := '0';
    P27RO2	: out std_logic := '0';
    P27RO3	: out std_logic := '0';
    P27RO4	: out std_logic := '0';
    P27RO5	: out std_logic := '0';

    P28CI1	: in std_logic := '0';
    P28CL	: in std_logic := '0';
    P28CR	: in std_logic := '0';
    P28CO	: out std_logic := '0';
    P28CTI	: in std_logic := '0';
    P28CTO	: out std_logic := '0';
    P28EI1	: in std_logic := '0';
    P28EI2	: in std_logic := '0';
    P28EI3	: in std_logic := '0';
    P28EI4	: in std_logic := '0';
    P28EI5	: in std_logic := '0';
    P28EL	: in std_logic := '0';
    P28ER	: in std_logic := '0';
    P28EO	: out std_logic := '0';
    P28RI	: in std_logic := '0';
    P28RL	: in std_logic := '0';
    P28RR	: in std_logic := '0';
    P28RO1	: out std_logic := '0';
    P28RO2	: out std_logic := '0';
    P28RO3	: out std_logic := '0';
    P28RO4	: out std_logic := '0';
    P28RO5	: out std_logic := '0';

    P29CI1	: in std_logic := '0';
    P29CL	: in std_logic := '0';
    P29CR	: in std_logic := '0';
    P29CO	: out std_logic := '0';
    P29CTI	: in std_logic := '0';
    P29CTO	: out std_logic := '0';
    P29EI1	: in std_logic := '0';
    P29EI2	: in std_logic := '0';
    P29EI3	: in std_logic := '0';
    P29EI4	: in std_logic := '0';
    P29EI5	: in std_logic := '0';
    P29EL	: in std_logic := '0';
    P29ER	: in std_logic := '0';
    P29EO	: out std_logic := '0';
    P29RI	: in std_logic := '0';
    P29RL	: in std_logic := '0';
    P29RR	: in std_logic := '0';
    P29RO1	: out std_logic := '0';
    P29RO2	: out std_logic := '0';
    P29RO3	: out std_logic := '0';
    P29RO4	: out std_logic := '0';
    P29RO5	: out std_logic := '0';

    P30CI1	: in std_logic := '0';
    P30CL	: in std_logic := '0';
    P30CR	: in std_logic := '0';
    P30CO	: out std_logic := '0';
    P30CTI	: in std_logic := '0';
    P30CTO	: out std_logic := '0';
    P30EI1	: in std_logic := '0';
    P30EI2	: in std_logic := '0';
    P30EI3	: in std_logic := '0';
    P30EI4	: in std_logic := '0';
    P30EI5	: in std_logic := '0';
    P30EL	: in std_logic := '0';
    P30ER	: in std_logic := '0';
    P30EO	: out std_logic := '0';
    P30RI	: in std_logic := '0';
    P30RL	: in std_logic := '0';
    P30RR	: in std_logic := '0';
    P30RO1	: out std_logic := '0';
    P30RO2	: out std_logic := '0';
    P30RO3	: out std_logic := '0';
    P30RO4	: out std_logic := '0';
    P30RO5	: out std_logic := '0'
);
end component NX_IOM;

component NX_IOM_CONTROL_M is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port (
    RTCK1	: in std_logic := '0';
    RRCK1	: in std_logic := '0';
    WTCK1	: in std_logic := '0';
    WRCK1	: in std_logic := '0';
    RTCK2	: in std_logic := '0';
    RRCK2	: in std_logic := '0';
    WTCK2	: in std_logic := '0';
    WRCK2	: in std_logic := '0';
    CTCK	: in std_logic := '0';

    C1TW	: in std_logic := '0';
    C1TS	: in std_logic := '0';
    C1RW1	: in std_logic := '0';
    C1RW2	: in std_logic := '0';
    C1RW3	: in std_logic := '0';
    C1RNE	: in std_logic := '0';
    C1RS	: in std_logic := '0';
    C2TW	: in std_logic := '0';
    C2TS	: in std_logic := '0';
    C2RW1	: in std_logic := '0';
    C2RW2	: in std_logic := '0';
    C2RW3	: in std_logic := '0';
    C2RNE	: in std_logic := '0';
    C2RS	: in std_logic := '0';
    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';
    DC	: in std_logic := '0';
    CCK	: in std_logic := '0';
    DCK	: in std_logic := '0';
    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';
    DRA5	: in std_logic := '0';
    DRA6	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DOS	: in std_logic := '0';
    DOG	: in std_logic := '0';
    DIS	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DPAS	: in std_logic := '0';
    DPAG	: in std_logic := '0';
    DQSS	: in std_logic := '0';
    DQSG	: in std_logic := '0';
    DS1	: in std_logic := '0';
    DS2	: in std_logic := '0';
    CAD1	: in std_logic := '0';
    CAD2	: in std_logic := '0';
    CAD3	: in std_logic := '0';
    CAD4	: in std_logic := '0';
    CAD5	: in std_logic := '0';
    CAD6	: in std_logic := '0';
    CAP1	: in std_logic := '0';
    CAP2	: in std_logic := '0';
    CAP3	: in std_logic := '0';
    CAP4	: in std_logic := '0';
    CAN1	: in std_logic := '0';
    CAN2	: in std_logic := '0';
    CAN3	: in std_logic := '0';
    CAN4	: in std_logic := '0';
    CAT1	: in std_logic := '0';
    CAT2	: in std_logic := '0';
    CAT3	: in std_logic := '0';
    CAT4	: in std_logic := '0';
    SPI1	: in std_logic := '0';
    SPI2	: in std_logic := '0';
    SPI3	: in std_logic := '0';
    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    C1RED	: out std_logic := '0';
    C2RED	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';
    CAL	: out std_logic := '0';

    LINK1	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK2	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK3	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK4	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK5	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK6	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK7	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK8	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK9	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK10	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK11	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK12	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK13	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK14	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK15	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK16	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK17	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK18	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK19	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK20	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK21	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK22	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK23	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK24	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK25	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK26	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK27	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK28	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK29	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK30	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK31	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK32	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK33	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK34	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_CONTROL_M;

component NX_IOM_DRIVER_U is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_type      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_type      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_type      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit := '0';

    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1	: in std_logic := '0';
    EI2	: in std_logic := '0';
    EI3	: in std_logic := '0';
    EI4	: in std_logic := '0';
    EI5	: in std_logic := '0';
    EI6	: in std_logic := '0';
    EI7	: in std_logic := '0';
    EI8	: in std_logic := '0';
    EL	: in std_logic := '0';
    ER	: in std_logic := '0';
    CI1	: in std_logic := '0';
    CL	: in std_logic := '0';
    CR	: in std_logic := '0';
    RI	: in std_logic := '0';
    RL	: in std_logic := '0';
    RR	: in std_logic := '0';
    CO	: out std_logic := '0';
    CTI	: in std_logic := '0';
    CTO	: out std_logic := '0';
    EO	: out std_logic := '0';
    RO1	: out std_logic := '0';
    RO2	: out std_logic := '0';
    RO3	: out std_logic := '0';
    RO4	: out std_logic := '0';
    RO5	: out std_logic := '0';
    RO6	: out std_logic := '0';
    RO7	: out std_logic := '0';
    RO8	: out std_logic := '0';
    LINK	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_DRIVER_U;

component NX_IOM_BIN2GRP is
port (
    LA	: in std_logic_vector(5 downto 0) := (others => '0');
    DS	: in std_logic_vector(1 downto 0) := (others => '0');

    GS	: in std_logic := '0';

    GVON	: out std_logic_vector(2 downto 0) := (others => '0');
    GVIN	: out std_logic_vector(2 downto 0) := (others => '0');
    GVDN	: out std_logic_vector(2 downto 0) := (others => '0');
    PA	: out std_logic_vector(3 downto 0) := (others => '0')
);
end component NX_IOM_BIN2GRP;

component NX_IOM_SERDES_U is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    FCK	: in std_logic := '0';
    SCK	: in std_logic := '0';
    LDRN	: in std_logic := '0';

    DRWDS	: in std_logic := '0';
    DRWEN	: in std_logic := '0';
    DRE	: in std_logic := '0';
    DRON	: in std_logic_vector(2 downto 0) := (others => '0');
    DRIN	: in std_logic_vector(2 downto 0) := (others => '0');
    DRDN	: in std_logic_vector(2 downto 0) := (others => '0');
    DRA	: in std_logic_vector(3 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');

    FA	: in std_logic_vector(5 downto 0) := (others => '0');
    FZ	: in std_logic := '0';

    ALD	: out std_logic := '0';
    ALT	: out std_logic := '0';

    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0');

    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';

    LINK	: inout std_logic_vector(IOM_LINK_SIZE-1 downto 0) := (others => '0')
);
end component NX_IOM_SERDES_U;

component NX_IOM_U is
generic (
    mode_side1        : integer := 0;
    div1         : bit_vector(2 downto 0) := "000";
    mode_side2        : integer := 0;
    div2         : bit_vector(2 downto 0) := "000";
    mode_side3        : integer := 0;
    div3         : bit_vector(2 downto 0) := "000";

    div_swrx1    : bit_vector(2 downto 0) := "000";
    div_swrx2    : bit_vector(2 downto 0) := "000";

    sel_ld_fck1  : bit_vector(1 downto 0) := "00";
    sel_ld_fck2  : bit_vector(1 downto 0) := "00";
    sel_ld_fck3  : bit_vector(1 downto 0) := "00";
    sel_sw_fck1  : bit_vector(1 downto 0) := "00";
    sel_sw_fck2  : bit_vector(1 downto 0) := "00";

    sel_dc_clk   : bit_vector(1 downto 0) := "00";

    inv_ld_sck1  : bit := '0';
    inv_ld_sck2  : bit := '0';
    inv_ld_sck3  : bit := '0';

    link_ld_12   : bit := '0';
    link_ld_23   : bit := '0';

    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';

    use_dc       : bit := '0';
    cal_delay1   : string := "";
    cal_delay2   : string := "";

    pads_dict    : string := "";
    pads_path    : string := ""
);
port (
    ALCK1	: in std_logic := '0';
    ALCK2	: in std_logic := '0';
    ALCK3	: in std_logic := '0';
    LDSCK1	: in std_logic := '0';
    LDSCK2	: in std_logic := '0';
    LDSCK3	: in std_logic := '0';
--  LDFCK1  : in    std_logic;	-- CONFIG
--  LDFCK2  : in    std_logic;	-- CONFIG
--  LDFCK3  : in    std_logic;	-- CONFIG
--  SWTX1CK : in    std_logic;	-- CONFIG
--  SWTX2CK : in    std_logic;	-- CONFIG
    SWRX1CK	: in std_logic := '0';
    SWRX2CK	: in std_logic := '0';
    FCK1	: in std_logic := '0';
    FCK2	: in std_logic := '0';
    FDCK	: in std_logic := '0';
    CCK	: in std_logic := '0';

    DQ1CI1	: in std_logic := '0';
    DQ1CI2	: in std_logic := '0';
    DQ1CI3	: in std_logic := '0';
    DQ1CI4	: in std_logic := '0';
    DQ1CI5	: in std_logic := '0';
    DQ1CI6	: in std_logic := '0';
    DQ1CI7	: in std_logic := '0';
    DQ1CI8	: in std_logic := '0';
    DQ2CI1	: in std_logic := '0';
    DQ2CI2	: in std_logic := '0';
    DQ2CI3	: in std_logic := '0';
    DQ2CI4	: in std_logic := '0';
    DQ2CI5	: in std_logic := '0';
    DQ2CI6	: in std_logic := '0';
    DQ2CI7	: in std_logic := '0';
    DQ2CI8	: in std_logic := '0';
    DQ3CI1	: in std_logic := '0';
    DQ3CI2	: in std_logic := '0';
    DQ3CI3	: in std_logic := '0';
    DQ3CI4	: in std_logic := '0';
    DQ3CI5	: in std_logic := '0';
    DQ3CI6	: in std_logic := '0';
    DQ3CI7	: in std_logic := '0';
    DQ3CI8	: in std_logic := '0';
    DQS1CI1	: in std_logic := '0';
    DQS1CI2	: in std_logic := '0';
    DQS1CI3	: in std_logic := '0';
    DQS1CI4	: in std_logic := '0';
    DQS1CI5	: in std_logic := '0';
    DQS1CI6	: in std_logic := '0';
    DQS1CI7	: in std_logic := '0';
    DQS1CI8	: in std_logic := '0';
    DQS2CI1	: in std_logic := '0';
    DQS2CI2	: in std_logic := '0';
    DQS2CI3	: in std_logic := '0';
    DQS2CI4	: in std_logic := '0';
    DQS2CI5	: in std_logic := '0';
    DQS2CI6	: in std_logic := '0';
    DQS2CI7	: in std_logic := '0';
    DQS2CI8	: in std_logic := '0';
    DQS3CI1	: in std_logic := '0';
    DQS3CI2	: in std_logic := '0';
    DQS3CI3	: in std_logic := '0';
    DQS3CI4	: in std_logic := '0';
    DQS3CI5	: in std_logic := '0';
    DQS3CI6	: in std_logic := '0';
    DQS3CI7	: in std_logic := '0';
    DQS3CI8	: in std_logic := '0';

    LD1RN	: in std_logic := '0';
    LD2RN	: in std_logic := '0';
    LD3RN	: in std_logic := '0';

    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';

    DCRN	: in std_logic := '0';
    LE	: in std_logic := '0';
    SE	: in std_logic := '0';

    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';

    DRO1CSN	: in std_logic := '0';
    DRO2CSN	: in std_logic := '0';
    DRO3CSN	: in std_logic := '0';
    DRI1CSN	: in std_logic := '0';
    DRI2CSN	: in std_logic := '0';
    DRI3CSN	: in std_logic := '0';
    DRDPA1CSN	: in std_logic := '0';
    DRDPA2CSN	: in std_logic := '0';
    DRDPA3CSN	: in std_logic := '0';
    DRCCSN	: in std_logic := '0';
    DRWDS	: in std_logic := '0';
    DRWEN	: in std_logic := '0';
    DRE	: in std_logic := '0';

    CA1P1	: in std_logic := '0';
    CA1P2	: in std_logic := '0';
    CA1P3	: in std_logic := '0';
    CA1P4	: in std_logic := '0';
    CA2P1	: in std_logic := '0';
    CA2P2	: in std_logic := '0';
    CA2P3	: in std_logic := '0';
    CA2P4	: in std_logic := '0';
    CA1N1	: in std_logic := '0';
    CA1N2	: in std_logic := '0';
    CA1N3	: in std_logic := '0';
    CA1N4	: in std_logic := '0';
    CA2N1	: in std_logic := '0';
    CA2N2	: in std_logic := '0';
    CA2N3	: in std_logic := '0';
    CA2N4	: in std_logic := '0';
    CA1T1	: in std_logic := '0';
    CA1T2	: in std_logic := '0';
    CA1T3	: in std_logic := '0';
    CA1T4	: in std_logic := '0';
    CA2T1	: in std_logic := '0';
    CA2T2	: in std_logic := '0';
    CA2T3	: in std_logic := '0';
    CA2T4	: in std_logic := '0';
    CA1D1	: in std_logic := '0';
    CA1D2	: in std_logic := '0';
    CA1D3	: in std_logic := '0';
    CA1D4	: in std_logic := '0';
    CA1D5	: in std_logic := '0';
    CA1D6	: in std_logic := '0';
    CA2D1	: in std_logic := '0';
    CA2D2	: in std_logic := '0';
    CA2D3	: in std_logic := '0';
    CA2D4	: in std_logic := '0';
    CA2D5	: in std_logic := '0';
    CA2D6	: in std_logic := '0';

    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';

    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    AL1D	: out std_logic := '0';
    AL2D	: out std_logic := '0';
    AL3D	: out std_logic := '0';
    AL1T	: out std_logic := '0';
    AL2T	: out std_logic := '0';
    AL3T	: out std_logic := '0';
    DCL	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';

    P1CI1	: in std_logic := '0';
    P1CL	: in std_logic := '0';
    P1CR	: in std_logic := '0';
    P1CO	: out std_logic := '0';
    P1CTI	: in std_logic := '0';
    P1CTO	: out std_logic := '0';
    P1EI1	: in std_logic := '0';
    P1EI2	: in std_logic := '0';
    P1EI3	: in std_logic := '0';
    P1EI4	: in std_logic := '0';
    P1EI5	: in std_logic := '0';
    P1EI6	: in std_logic := '0';
    P1EI7	: in std_logic := '0';
    P1EI8	: in std_logic := '0';

    P1EL	: in std_logic := '0';
    P1ER	: in std_logic := '0';
    P1EO	: out std_logic := '0';
    P1RI	: in std_logic := '0';
    P1RL	: in std_logic := '0';
    P1RR	: in std_logic := '0';
    P1RO1	: out std_logic := '0';
    P1RO2	: out std_logic := '0';
    P1RO3	: out std_logic := '0';
    P1RO4	: out std_logic := '0';
    P1RO5	: out std_logic := '0';
    P1RO6	: out std_logic := '0';
    P1RO7	: out std_logic := '0';
    P1RO8	: out std_logic := '0';

    P2CI1	: in std_logic := '0';
    P2CL	: in std_logic := '0';
    P2CR	: in std_logic := '0';
    P2CO	: out std_logic := '0';
    P2CTI	: in std_logic := '0';
    P2CTO	: out std_logic := '0';
    P2EI1	: in std_logic := '0';
    P2EI2	: in std_logic := '0';
    P2EI3	: in std_logic := '0';
    P2EI4	: in std_logic := '0';
    P2EI5	: in std_logic := '0';
    P2EI6	: in std_logic := '0';
    P2EI7	: in std_logic := '0';
    P2EI8	: in std_logic := '0';

    P2EL	: in std_logic := '0';
    P2ER	: in std_logic := '0';
    P2EO	: out std_logic := '0';
    P2RI	: in std_logic := '0';
    P2RL	: in std_logic := '0';
    P2RR	: in std_logic := '0';
    P2RO1	: out std_logic := '0';
    P2RO2	: out std_logic := '0';
    P2RO3	: out std_logic := '0';
    P2RO4	: out std_logic := '0';
    P2RO5	: out std_logic := '0';
    P2RO6	: out std_logic := '0';
    P2RO7	: out std_logic := '0';
    P2RO8	: out std_logic := '0';

    P3CI1	: in std_logic := '0';
    P3CL	: in std_logic := '0';
    P3CR	: in std_logic := '0';
    P3CO	: out std_logic := '0';
    P3CTI	: in std_logic := '0';
    P3CTO	: out std_logic := '0';
    P3EI1	: in std_logic := '0';
    P3EI2	: in std_logic := '0';
    P3EI3	: in std_logic := '0';
    P3EI4	: in std_logic := '0';
    P3EI5	: in std_logic := '0';
    P3EI6	: in std_logic := '0';
    P3EI7	: in std_logic := '0';
    P3EI8	: in std_logic := '0';

    P3EL	: in std_logic := '0';
    P3ER	: in std_logic := '0';
    P3EO	: out std_logic := '0';
    P3RI	: in std_logic := '0';
    P3RL	: in std_logic := '0';
    P3RR	: in std_logic := '0';
    P3RO1	: out std_logic := '0';
    P3RO2	: out std_logic := '0';
    P3RO3	: out std_logic := '0';
    P3RO4	: out std_logic := '0';
    P3RO5	: out std_logic := '0';
    P3RO6	: out std_logic := '0';
    P3RO7	: out std_logic := '0';
    P3RO8	: out std_logic := '0';

    P4CI1	: in std_logic := '0';
    P4CL	: in std_logic := '0';
    P4CR	: in std_logic := '0';
    P4CO	: out std_logic := '0';
    P4CTI	: in std_logic := '0';
    P4CTO	: out std_logic := '0';
    P4EI1	: in std_logic := '0';
    P4EI2	: in std_logic := '0';
    P4EI3	: in std_logic := '0';
    P4EI4	: in std_logic := '0';
    P4EI5	: in std_logic := '0';
    P4EI6	: in std_logic := '0';
    P4EI7	: in std_logic := '0';
    P4EI8	: in std_logic := '0';

    P4EL	: in std_logic := '0';
    P4ER	: in std_logic := '0';
    P4EO	: out std_logic := '0';
    P4RI	: in std_logic := '0';
    P4RL	: in std_logic := '0';
    P4RR	: in std_logic := '0';
    P4RO1	: out std_logic := '0';
    P4RO2	: out std_logic := '0';
    P4RO3	: out std_logic := '0';
    P4RO4	: out std_logic := '0';
    P4RO5	: out std_logic := '0';
    P4RO6	: out std_logic := '0';
    P4RO7	: out std_logic := '0';
    P4RO8	: out std_logic := '0';

    P5CI1	: in std_logic := '0';
    P5CL	: in std_logic := '0';
    P5CR	: in std_logic := '0';
    P5CO	: out std_logic := '0';
    P5CTI	: in std_logic := '0';
    P5CTO	: out std_logic := '0';
    P5EI1	: in std_logic := '0';
    P5EI2	: in std_logic := '0';
    P5EI3	: in std_logic := '0';
    P5EI4	: in std_logic := '0';
    P5EI5	: in std_logic := '0';
    P5EI6	: in std_logic := '0';
    P5EI7	: in std_logic := '0';
    P5EI8	: in std_logic := '0';

    P5EL	: in std_logic := '0';
    P5ER	: in std_logic := '0';
    P5EO	: out std_logic := '0';
    P5RI	: in std_logic := '0';
    P5RL	: in std_logic := '0';
    P5RR	: in std_logic := '0';
    P5RO1	: out std_logic := '0';
    P5RO2	: out std_logic := '0';
    P5RO3	: out std_logic := '0';
    P5RO4	: out std_logic := '0';
    P5RO5	: out std_logic := '0';
    P5RO6	: out std_logic := '0';
    P5RO7	: out std_logic := '0';
    P5RO8	: out std_logic := '0';

    P6CI1	: in std_logic := '0';
    P6CL	: in std_logic := '0';
    P6CR	: in std_logic := '0';
    P6CO	: out std_logic := '0';
    P6CTI	: in std_logic := '0';
    P6CTO	: out std_logic := '0';
    P6EI1	: in std_logic := '0';
    P6EI2	: in std_logic := '0';
    P6EI3	: in std_logic := '0';
    P6EI4	: in std_logic := '0';
    P6EI5	: in std_logic := '0';
    P6EI6	: in std_logic := '0';
    P6EI7	: in std_logic := '0';
    P6EI8	: in std_logic := '0';

    P6EL	: in std_logic := '0';
    P6ER	: in std_logic := '0';
    P6EO	: out std_logic := '0';
    P6RI	: in std_logic := '0';
    P6RL	: in std_logic := '0';
    P6RR	: in std_logic := '0';
    P6RO1	: out std_logic := '0';
    P6RO2	: out std_logic := '0';
    P6RO3	: out std_logic := '0';
    P6RO4	: out std_logic := '0';
    P6RO5	: out std_logic := '0';
    P6RO6	: out std_logic := '0';
    P6RO7	: out std_logic := '0';
    P6RO8	: out std_logic := '0';

    P7CI1	: in std_logic := '0';
    P7CL	: in std_logic := '0';
    P7CR	: in std_logic := '0';
    P7CO	: out std_logic := '0';
    P7CTI	: in std_logic := '0';
    P7CTO	: out std_logic := '0';
    P7EI1	: in std_logic := '0';
    P7EI2	: in std_logic := '0';
    P7EI3	: in std_logic := '0';
    P7EI4	: in std_logic := '0';
    P7EI5	: in std_logic := '0';
    P7EI6	: in std_logic := '0';
    P7EI7	: in std_logic := '0';
    P7EI8	: in std_logic := '0';

    P7EL	: in std_logic := '0';
    P7ER	: in std_logic := '0';
    P7EO	: out std_logic := '0';
    P7RI	: in std_logic := '0';
    P7RL	: in std_logic := '0';
    P7RR	: in std_logic := '0';
    P7RO1	: out std_logic := '0';
    P7RO2	: out std_logic := '0';
    P7RO3	: out std_logic := '0';
    P7RO4	: out std_logic := '0';
    P7RO5	: out std_logic := '0';
    P7RO6	: out std_logic := '0';
    P7RO7	: out std_logic := '0';
    P7RO8	: out std_logic := '0';

    P8CI1	: in std_logic := '0';
    P8CL	: in std_logic := '0';
    P8CR	: in std_logic := '0';
    P8CO	: out std_logic := '0';
    P8CTI	: in std_logic := '0';
    P8CTO	: out std_logic := '0';
    P8EI1	: in std_logic := '0';
    P8EI2	: in std_logic := '0';
    P8EI3	: in std_logic := '0';
    P8EI4	: in std_logic := '0';
    P8EI5	: in std_logic := '0';
    P8EI6	: in std_logic := '0';
    P8EI7	: in std_logic := '0';
    P8EI8	: in std_logic := '0';

    P8EL	: in std_logic := '0';
    P8ER	: in std_logic := '0';
    P8EO	: out std_logic := '0';
    P8RI	: in std_logic := '0';
    P8RL	: in std_logic := '0';
    P8RR	: in std_logic := '0';
    P8RO1	: out std_logic := '0';
    P8RO2	: out std_logic := '0';
    P8RO3	: out std_logic := '0';
    P8RO4	: out std_logic := '0';
    P8RO5	: out std_logic := '0';
    P8RO6	: out std_logic := '0';
    P8RO7	: out std_logic := '0';
    P8RO8	: out std_logic := '0';

    P9CI1	: in std_logic := '0';
    P9CL	: in std_logic := '0';
    P9CR	: in std_logic := '0';
    P9CO	: out std_logic := '0';
    P9CTI	: in std_logic := '0';
    P9CTO	: out std_logic := '0';
    P9EI1	: in std_logic := '0';
    P9EI2	: in std_logic := '0';
    P9EI3	: in std_logic := '0';
    P9EI4	: in std_logic := '0';
    P9EI5	: in std_logic := '0';
    P9EI6	: in std_logic := '0';
    P9EI7	: in std_logic := '0';
    P9EI8	: in std_logic := '0';

    P9EL	: in std_logic := '0';
    P9ER	: in std_logic := '0';
    P9EO	: out std_logic := '0';
    P9RI	: in std_logic := '0';
    P9RL	: in std_logic := '0';
    P9RR	: in std_logic := '0';
    P9RO1	: out std_logic := '0';
    P9RO2	: out std_logic := '0';
    P9RO3	: out std_logic := '0';
    P9RO4	: out std_logic := '0';
    P9RO5	: out std_logic := '0';
    P9RO6	: out std_logic := '0';
    P9RO7	: out std_logic := '0';
    P9RO8	: out std_logic := '0';

    P10CI1	: in std_logic := '0';
    P10CL	: in std_logic := '0';
    P10CR	: in std_logic := '0';
    P10CO	: out std_logic := '0';
    P10CTI	: in std_logic := '0';
    P10CTO	: out std_logic := '0';
    P10EI1	: in std_logic := '0';
    P10EI2	: in std_logic := '0';
    P10EI3	: in std_logic := '0';
    P10EI4	: in std_logic := '0';
    P10EI5	: in std_logic := '0';
    P10EI6	: in std_logic := '0';
    P10EI7	: in std_logic := '0';
    P10EI8	: in std_logic := '0';

    P10EL	: in std_logic := '0';
    P10ER	: in std_logic := '0';
    P10EO	: out std_logic := '0';
    P10RI	: in std_logic := '0';
    P10RL	: in std_logic := '0';
    P10RR	: in std_logic := '0';
    P10RO1	: out std_logic := '0';
    P10RO2	: out std_logic := '0';
    P10RO3	: out std_logic := '0';
    P10RO4	: out std_logic := '0';
    P10RO5	: out std_logic := '0';
    P10RO6	: out std_logic := '0';
    P10RO7	: out std_logic := '0';
    P10RO8	: out std_logic := '0';

    P11CI1	: in std_logic := '0';
    
    P11CL	: in std_logic := '0';
    P11CR	: in std_logic := '0';
    P11CO	: out std_logic := '0';
    P11CTI	: in std_logic := '0';
    P11CTO	: out std_logic := '0';
    P11EI1	: in std_logic := '0';
    P11EI2	: in std_logic := '0';
    P11EI3	: in std_logic := '0';
    P11EI4	: in std_logic := '0';
    P11EI5	: in std_logic := '0';
    P11EI6	: in std_logic := '0';
    P11EI7	: in std_logic := '0';
    P11EI8	: in std_logic := '0';

    P11EL	: in std_logic := '0';
    P11ER	: in std_logic := '0';
    P11EO	: out std_logic := '0';
    P11RI	: in std_logic := '0';
    P11RL	: in std_logic := '0';
    P11RR	: in std_logic := '0';
    P11RO1	: out std_logic := '0';
    P11RO2	: out std_logic := '0';
    P11RO3	: out std_logic := '0';
    P11RO4	: out std_logic := '0';
    P11RO5	: out std_logic := '0';
    P11RO6	: out std_logic := '0';
    P11RO7	: out std_logic := '0';
    P11RO8	: out std_logic := '0';

    P12CI1	: in std_logic := '0';
    P12CL	: in std_logic := '0';
    P12CR	: in std_logic := '0';
    P12CO	: out std_logic := '0';
    P12CTI	: in std_logic := '0';
    P12CTO	: out std_logic := '0';
    P12EI1	: in std_logic := '0';
    P12EI2	: in std_logic := '0';
    P12EI3	: in std_logic := '0';
    P12EI4	: in std_logic := '0';
    P12EI5	: in std_logic := '0';
    P12EI6	: in std_logic := '0';
    P12EI7	: in std_logic := '0';
    P12EI8	: in std_logic := '0';

    P12EL	: in std_logic := '0';
    P12ER	: in std_logic := '0';
    P12EO	: out std_logic := '0';
    P12RI	: in std_logic := '0';
    P12RL	: in std_logic := '0';
    P12RR	: in std_logic := '0';
    P12RO1	: out std_logic := '0';
    P12RO2	: out std_logic := '0';
    P12RO3	: out std_logic := '0';
    P12RO4	: out std_logic := '0';
    P12RO5	: out std_logic := '0';
    P12RO6	: out std_logic := '0';
    P12RO7	: out std_logic := '0';
    P12RO8	: out std_logic := '0';

    P13CI1	: in std_logic := '0';
    P13CL	: in std_logic := '0';
    P13CR	: in std_logic := '0';
    P13CO	: out std_logic := '0';
    P13CTI	: in std_logic := '0';
    P13CTO	: out std_logic := '0';
    P13EI1	: in std_logic := '0';
    P13EI2	: in std_logic := '0';
    P13EI3	: in std_logic := '0';
    P13EI4	: in std_logic := '0';
    P13EI5	: in std_logic := '0';
    P13EI6	: in std_logic := '0';
    P13EI7	: in std_logic := '0';
    P13EI8	: in std_logic := '0';

    P13EL	: in std_logic := '0';
    P13ER	: in std_logic := '0';
    P13EO	: out std_logic := '0';
    P13RI	: in std_logic := '0';
    P13RL	: in std_logic := '0';
    P13RR	: in std_logic := '0';
    P13RO1	: out std_logic := '0';
    P13RO2	: out std_logic := '0';
    P13RO3	: out std_logic := '0';
    P13RO4	: out std_logic := '0';
    P13RO5	: out std_logic := '0';
    P13RO6	: out std_logic := '0';
    P13RO7	: out std_logic := '0';
    P13RO8	: out std_logic := '0';

    P14CI1	: in std_logic := '0';
    P14CL	: in std_logic := '0';
    P14CR	: in std_logic := '0';
    P14CO	: out std_logic := '0';
    P14CTI	: in std_logic := '0';
    P14CTO	: out std_logic := '0';
    P14EI1	: in std_logic := '0';
    P14EI2	: in std_logic := '0';
    P14EI3	: in std_logic := '0';
    P14EI4	: in std_logic := '0';
    P14EI5	: in std_logic := '0';
    P14EI6	: in std_logic := '0';
    P14EI7	: in std_logic := '0';
    P14EI8	: in std_logic := '0';

    P14EL	: in std_logic := '0';
    P14ER	: in std_logic := '0';
    P14EO	: out std_logic := '0';
    P14RI	: in std_logic := '0';
    P14RL	: in std_logic := '0';
    P14RR	: in std_logic := '0';
    P14RO1	: out std_logic := '0';
    P14RO2	: out std_logic := '0';
    P14RO3	: out std_logic := '0';
    P14RO4	: out std_logic := '0';
    P14RO5	: out std_logic := '0';
    P14RO6	: out std_logic := '0';
    P14RO7	: out std_logic := '0';
    P14RO8	: out std_logic := '0';

    P15CI1	: in std_logic := '0';
    P15CL	: in std_logic := '0';
    P15CR	: in std_logic := '0';
    P15CO	: out std_logic := '0';
    P15CTI	: in std_logic := '0';
    P15CTO	: out std_logic := '0';
    P15EI1	: in std_logic := '0';
    P15EI2	: in std_logic := '0';
    P15EI3	: in std_logic := '0';
    P15EI4	: in std_logic := '0';
    P15EI5	: in std_logic := '0';
    P15EI6	: in std_logic := '0';
    P15EI7	: in std_logic := '0';
    P15EI8	: in std_logic := '0';

    P15EL	: in std_logic := '0';
    P15ER	: in std_logic := '0';
    P15EO	: out std_logic := '0';
    P15RI	: in std_logic := '0';
    P15RL	: in std_logic := '0';
    P15RR	: in std_logic := '0';
    P15RO1	: out std_logic := '0';
    P15RO2	: out std_logic := '0';
    P15RO3	: out std_logic := '0';
    P15RO4	: out std_logic := '0';
    P15RO5	: out std_logic := '0';
    P15RO6	: out std_logic := '0';
    P15RO7	: out std_logic := '0';
    P15RO8	: out std_logic := '0';

    P16CI1	: in std_logic := '0';
    P16CL	: in std_logic := '0';
    P16CR	: in std_logic := '0';
    P16CO	: out std_logic := '0';
    P16CTI	: in std_logic := '0';
    P16CTO	: out std_logic := '0';
    P16EI1	: in std_logic := '0';
    P16EI2	: in std_logic := '0';
    P16EI3	: in std_logic := '0';
    P16EI4	: in std_logic := '0';
    P16EI5	: in std_logic := '0';
    P16EI6	: in std_logic := '0';
    P16EI7	: in std_logic := '0';
    P16EI8	: in std_logic := '0';

    P16EL	: in std_logic := '0';
    P16ER	: in std_logic := '0';
    P16EO	: out std_logic := '0';
    P16RI	: in std_logic := '0';
    P16RL	: in std_logic := '0';
    P16RR	: in std_logic := '0';
    P16RO1	: out std_logic := '0';
    P16RO2	: out std_logic := '0';
    P16RO3	: out std_logic := '0';
    P16RO4	: out std_logic := '0';
    P16RO5	: out std_logic := '0';
    P16RO6	: out std_logic := '0';
    P16RO7	: out std_logic := '0';
    P16RO8	: out std_logic := '0';

    P17CI1	: in std_logic := '0';
    P17CL	: in std_logic := '0';
    P17CR	: in std_logic := '0';
    P17CO	: out std_logic := '0';
    P17CTI	: in std_logic := '0';
    P17CTO	: out std_logic := '0';
    P17EI1	: in std_logic := '0';
    P17EI2	: in std_logic := '0';
    P17EI3	: in std_logic := '0';
    P17EI4	: in std_logic := '0';
    P17EI5	: in std_logic := '0';
    P17EI6	: in std_logic := '0';
    P17EI7	: in std_logic := '0';
    P17EI8	: in std_logic := '0';

    P17EL	: in std_logic := '0';
    P17ER	: in std_logic := '0';
    P17EO	: out std_logic := '0';
    P17RI	: in std_logic := '0';
    P17RL	: in std_logic := '0';
    P17RR	: in std_logic := '0';
    P17RO1	: out std_logic := '0';
    P17RO2	: out std_logic := '0';
    P17RO3	: out std_logic := '0';
    P17RO4	: out std_logic := '0';
    P17RO5	: out std_logic := '0';
    P17RO6	: out std_logic := '0';
    P17RO7	: out std_logic := '0';
    P17RO8	: out std_logic := '0';

    P18CI1	: in std_logic := '0';
    P18CL	: in std_logic := '0';
    P18CR	: in std_logic := '0';
    P18CO	: out std_logic := '0';
    P18CTI	: in std_logic := '0';
    P18CTO	: out std_logic := '0';
    P18EI1	: in std_logic := '0';
    P18EI2	: in std_logic := '0';
    P18EI3	: in std_logic := '0';
    P18EI4	: in std_logic := '0';
    P18EI5	: in std_logic := '0';
    P18EI6	: in std_logic := '0';
    P18EI7	: in std_logic := '0';
    P18EI8	: in std_logic := '0';

    P18EL	: in std_logic := '0';
    P18ER	: in std_logic := '0';
    P18EO	: out std_logic := '0';
    P18RI	: in std_logic := '0';
    P18RL	: in std_logic := '0';
    P18RR	: in std_logic := '0';
    P18RO1	: out std_logic := '0';
    P18RO2	: out std_logic := '0';
    P18RO3	: out std_logic := '0';
    P18RO4	: out std_logic := '0';
    P18RO5	: out std_logic := '0';
    P18RO6	: out std_logic := '0';
    P18RO7	: out std_logic := '0';
    P18RO8	: out std_logic := '0';

    P19CI1	: in std_logic := '0';
    P19CL	: in std_logic := '0';
    P19CR	: in std_logic := '0';
    P19CO	: out std_logic := '0';
    P19CTI	: in std_logic := '0';
    P19CTO	: out std_logic := '0';
    P19EI1	: in std_logic := '0';
    P19EI2	: in std_logic := '0';
    P19EI3	: in std_logic := '0';
    P19EI4	: in std_logic := '0';
    P19EI5	: in std_logic := '0';
    P19EI6	: in std_logic := '0';
    P19EI7	: in std_logic := '0';
    P19EI8	: in std_logic := '0';

    P19EL	: in std_logic := '0';
    P19ER	: in std_logic := '0';
    P19EO	: out std_logic := '0';
    P19RI	: in std_logic := '0';
    P19RL	: in std_logic := '0';
    P19RR	: in std_logic := '0';
    P19RO1	: out std_logic := '0';
    P19RO2	: out std_logic := '0';
    P19RO3	: out std_logic := '0';
    P19RO4	: out std_logic := '0';
    P19RO5	: out std_logic := '0';
    P19RO6	: out std_logic := '0';
    P19RO7	: out std_logic := '0';
    P19RO8	: out std_logic := '0';

    P20CI1	: in std_logic := '0';
    P20CL	: in std_logic := '0';
    P20CR	: in std_logic := '0';
    P20CO	: out std_logic := '0';
    P20CTI	: in std_logic := '0';
    P20CTO	: out std_logic := '0';
    P20EI1	: in std_logic := '0';
    P20EI2	: in std_logic := '0';
    P20EI3	: in std_logic := '0';
    P20EI4	: in std_logic := '0';
    P20EI5	: in std_logic := '0';
    P20EI6	: in std_logic := '0';
    P20EI7	: in std_logic := '0';
    P20EI8	: in std_logic := '0';

    P20EL	: in std_logic := '0';
    P20ER	: in std_logic := '0';
    P20EO	: out std_logic := '0';
    P20RI	: in std_logic := '0';
    P20RL	: in std_logic := '0';
    P20RR	: in std_logic := '0';
    P20RO1	: out std_logic := '0';
    P20RO2	: out std_logic := '0';
    P20RO3	: out std_logic := '0';
    P20RO4	: out std_logic := '0';
    P20RO5	: out std_logic := '0';
    P20RO6	: out std_logic := '0';
    P20RO7	: out std_logic := '0';
    P20RO8	: out std_logic := '0';

    P21CI1	: in std_logic := '0';
    P21CL	: in std_logic := '0';
    P21CR	: in std_logic := '0';
    P21CO	: out std_logic := '0';
    P21CTI	: in std_logic := '0';
    P21CTO	: out std_logic := '0';
    P21EI1	: in std_logic := '0';
    P21EI2	: in std_logic := '0';
    P21EI3	: in std_logic := '0';
    P21EI4	: in std_logic := '0';
    P21EI5	: in std_logic := '0';
    P21EI6	: in std_logic := '0';
    P21EI7	: in std_logic := '0';
    P21EI8	: in std_logic := '0';

    P21EL	: in std_logic := '0';
    P21ER	: in std_logic := '0';
    P21EO	: out std_logic := '0';
    P21RI	: in std_logic := '0';
    P21RL	: in std_logic := '0';
    P21RR	: in std_logic := '0';
    P21RO1	: out std_logic := '0';
    P21RO2	: out std_logic := '0';
    P21RO3	: out std_logic := '0';
    P21RO4	: out std_logic := '0';
    P21RO5	: out std_logic := '0';
    P21RO6	: out std_logic := '0';
    P21RO7	: out std_logic := '0';
    P21RO8	: out std_logic := '0';

    P22CI1	: in std_logic := '0';
    P22CL	: in std_logic := '0';
    P22CR	: in std_logic := '0';
    P22CO	: out std_logic := '0';
    P22CTI	: in std_logic := '0';
    P22CTO	: out std_logic := '0';
    P22EI1	: in std_logic := '0';
    P22EI2	: in std_logic := '0';
    P22EI3	: in std_logic := '0';
    P22EI4	: in std_logic := '0';
    P22EI5	: in std_logic := '0';
    P22EI6	: in std_logic := '0';
    P22EI7	: in std_logic := '0';
    P22EI8	: in std_logic := '0';

    P22EL	: in std_logic := '0';
    P22ER	: in std_logic := '0';
    P22EO	: out std_logic := '0';
    P22RI	: in std_logic := '0';
    P22RL	: in std_logic := '0';
    P22RR	: in std_logic := '0';
    P22RO1	: out std_logic := '0';
    P22RO2	: out std_logic := '0';
    P22RO3	: out std_logic := '0';
    P22RO4	: out std_logic := '0';
    P22RO5	: out std_logic := '0';
    P22RO6	: out std_logic := '0';
    P22RO7	: out std_logic := '0';
    P22RO8	: out std_logic := '0';

    P23CI1	: in std_logic := '0';
    P23CL	: in std_logic := '0';
    P23CR	: in std_logic := '0';
    P23CO	: out std_logic := '0';
    P23CTI	: in std_logic := '0';
    P23CTO	: out std_logic := '0';
    P23EI1	: in std_logic := '0';
    P23EI2	: in std_logic := '0';
    P23EI3	: in std_logic := '0';
    P23EI4	: in std_logic := '0';
    P23EI5	: in std_logic := '0';
    P23EI6	: in std_logic := '0';
    P23EI7	: in std_logic := '0';
    P23EI8	: in std_logic := '0';

    P23EL	: in std_logic := '0';
    P23ER	: in std_logic := '0';
    P23EO	: out std_logic := '0';
    P23RI	: in std_logic := '0';
    P23RL	: in std_logic := '0';
    P23RR	: in std_logic := '0';
    P23RO1	: out std_logic := '0';
    P23RO2	: out std_logic := '0';
    P23RO3	: out std_logic := '0';
    P23RO4	: out std_logic := '0';
    P23RO5	: out std_logic := '0';
    P23RO6	: out std_logic := '0';
    P23RO7	: out std_logic := '0';
    P23RO8	: out std_logic := '0';

    P24CI1	: in std_logic := '0';
    P24CL	: in std_logic := '0';
    P24CR	: in std_logic := '0';
    P24CO	: out std_logic := '0';
    P24CTI	: in std_logic := '0';
    P24CTO	: out std_logic := '0';
    P24EI1	: in std_logic := '0';
    P24EI2	: in std_logic := '0';
    P24EI3	: in std_logic := '0';
    P24EI4	: in std_logic := '0';
    P24EI5	: in std_logic := '0';
    P24EI6	: in std_logic := '0';
    P24EI7	: in std_logic := '0';
    P24EI8	: in std_logic := '0';

    P24EL	: in std_logic := '0';
    P24ER	: in std_logic := '0';
    P24EO	: out std_logic := '0';
    P24RI	: in std_logic := '0';
    P24RL	: in std_logic := '0';
    P24RR	: in std_logic := '0';
    P24RO1	: out std_logic := '0';
    P24RO2	: out std_logic := '0';
    P24RO3	: out std_logic := '0';
    P24RO4	: out std_logic := '0';
    P24RO5	: out std_logic := '0';
    P24RO6	: out std_logic := '0';
    P24RO7	: out std_logic := '0';
    P24RO8	: out std_logic := '0';

    P25CI1	: in std_logic := '0';
    P25CL	: in std_logic := '0';
    P25CR	: in std_logic := '0';
    P25CO	: out std_logic := '0';
    P25CTI	: in std_logic := '0';
    P25CTO	: out std_logic := '0';
    P25EI1	: in std_logic := '0';
    P25EI2	: in std_logic := '0';
    P25EI3	: in std_logic := '0';
    P25EI4	: in std_logic := '0';
    P25EI5	: in std_logic := '0';
    P25EI6	: in std_logic := '0';
    P25EI7	: in std_logic := '0';
    P25EI8	: in std_logic := '0';

    P25EL	: in std_logic := '0';
    P25ER	: in std_logic := '0';
    P25EO	: out std_logic := '0';
    P25RI	: in std_logic := '0';
    P25RL	: in std_logic := '0';
    P25RR	: in std_logic := '0';
    P25RO1	: out std_logic := '0';
    P25RO2	: out std_logic := '0';
    P25RO3	: out std_logic := '0';
    P25RO4	: out std_logic := '0';
    P25RO5	: out std_logic := '0';
    P25RO6	: out std_logic := '0';
    P25RO7	: out std_logic := '0';
    P25RO8	: out std_logic := '0';

    P26CI1	: in std_logic := '0';
    P26CL	: in std_logic := '0';
    P26CR	: in std_logic := '0';
    P26CO	: out std_logic := '0';
    P26CTI	: in std_logic := '0';
    P26CTO	: out std_logic := '0';
    P26EI1	: in std_logic := '0';
    P26EI2	: in std_logic := '0';
    P26EI3	: in std_logic := '0';
    P26EI4	: in std_logic := '0';
    P26EI5	: in std_logic := '0';
    P26EI6	: in std_logic := '0';
    P26EI7	: in std_logic := '0';
    P26EI8	: in std_logic := '0';

    P26EL	: in std_logic := '0';
    P26ER	: in std_logic := '0';
    P26EO	: out std_logic := '0';
    P26RI	: in std_logic := '0';
    P26RL	: in std_logic := '0';
    P26RR	: in std_logic := '0';
    P26RO1	: out std_logic := '0';
    P26RO2	: out std_logic := '0';
    P26RO3	: out std_logic := '0';
    P26RO4	: out std_logic := '0';
    P26RO5	: out std_logic := '0';
    P26RO6	: out std_logic := '0';
    P26RO7	: out std_logic := '0';
    P26RO8	: out std_logic := '0';

    P27CI1	: in std_logic := '0';
    P27CL	: in std_logic := '0';
    P27CR	: in std_logic := '0';
    P27CO	: out std_logic := '0';
    P27CTI	: in std_logic := '0';
    P27CTO	: out std_logic := '0';
    P27EI1	: in std_logic := '0';
    P27EI2	: in std_logic := '0';
    P27EI3	: in std_logic := '0';
    P27EI4	: in std_logic := '0';
    P27EI5	: in std_logic := '0';
    P27EI6	: in std_logic := '0';
    P27EI7	: in std_logic := '0';
    P27EI8	: in std_logic := '0';

    P27EL	: in std_logic := '0';
    P27ER	: in std_logic := '0';
    P27EO	: out std_logic := '0';
    P27RI	: in std_logic := '0';
    P27RL	: in std_logic := '0';
    P27RR	: in std_logic := '0';
    P27RO1	: out std_logic := '0';
    P27RO2	: out std_logic := '0';
    P27RO3	: out std_logic := '0';
    P27RO4	: out std_logic := '0';
    P27RO5	: out std_logic := '0';
    P27RO6	: out std_logic := '0';
    P27RO7	: out std_logic := '0';
    P27RO8	: out std_logic := '0';

    P28CI1	: in std_logic := '0';
    P28CL	: in std_logic := '0';
    P28CR	: in std_logic := '0';
    P28CO	: out std_logic := '0';
    P28CTI	: in std_logic := '0';
    P28CTO	: out std_logic := '0';
    P28EI1	: in std_logic := '0';
    P28EI2	: in std_logic := '0';
    P28EI3	: in std_logic := '0';
    P28EI4	: in std_logic := '0';
    P28EI5	: in std_logic := '0';
    P28EI6	: in std_logic := '0';
    P28EI7	: in std_logic := '0';
    P28EI8	: in std_logic := '0';
    P28EL	: in std_logic := '0';
    P28ER	: in std_logic := '0';
    P28EO	: out std_logic := '0';
    P28RI	: in std_logic := '0';
    P28RL	: in std_logic := '0';
    P28RR	: in std_logic := '0';
    P28RO1	: out std_logic := '0';
    P28RO2	: out std_logic := '0';
    P28RO3	: out std_logic := '0';
    P28RO4	: out std_logic := '0';
    P28RO5	: out std_logic := '0';
    P28RO6	: out std_logic := '0';
    P28RO7	: out std_logic := '0';
    P28RO8	: out std_logic := '0';

    P29CI1	: in std_logic := '0';
    P29CL	: in std_logic := '0';
    P29CR	: in std_logic := '0';
    P29CO	: out std_logic := '0';
    P29CTI	: in std_logic := '0';
    P29CTO	: out std_logic := '0';
    P29EI1	: in std_logic := '0';
    P29EI2	: in std_logic := '0';
    P29EI3	: in std_logic := '0';
    P29EI4	: in std_logic := '0';
    P29EI5	: in std_logic := '0';
    P29EI6	: in std_logic := '0';
    P29EI7	: in std_logic := '0';
    P29EI8	: in std_logic := '0';
    P29EL	: in std_logic := '0';
    P29ER	: in std_logic := '0';
    P29EO	: out std_logic := '0';
    P29RI	: in std_logic := '0';
    P29RL	: in std_logic := '0';
    P29RR	: in std_logic := '0';
    P29RO1	: out std_logic := '0';
    P29RO2	: out std_logic := '0';
    P29RO3	: out std_logic := '0';
    P29RO4	: out std_logic := '0';
    P29RO5	: out std_logic := '0';
    P29RO6	: out std_logic := '0';
    P29RO7	: out std_logic := '0';
    P29RO8	: out std_logic := '0';

    P30CI1	: in std_logic := '0';
    P30CL	: in std_logic := '0';
    P30CR	: in std_logic := '0';
    P30CO	: out std_logic := '0';
    P30CTI	: in std_logic := '0';
    P30CTO	: out std_logic := '0';
    P30EI1	: in std_logic := '0';
    P30EI2	: in std_logic := '0';
    P30EI3	: in std_logic := '0';
    P30EI4	: in std_logic := '0';
    P30EI5	: in std_logic := '0';
    P30EI6	: in std_logic := '0';
    P30EI7	: in std_logic := '0';
    P30EI8	: in std_logic := '0';
    P30EL	: in std_logic := '0';
    P30ER	: in std_logic := '0';
    P30EO	: out std_logic := '0';
    P30RI	: in std_logic := '0';
    P30RL	: in std_logic := '0';
    P30RR	: in std_logic := '0';
    P30RO1	: out std_logic := '0';
    P30RO2	: out std_logic := '0';
    P30RO3	: out std_logic := '0';
    P30RO4	: out std_logic := '0';
    P30RO5	: out std_logic := '0';
    P30RO6	: out std_logic := '0';
    P30RO7	: out std_logic := '0';
    P30RO8	: out std_logic := '0';

    P31CI1	: in std_logic := '0';
    P31CL	: in std_logic := '0';
    P31CR	: in std_logic := '0';
    P31CO	: out std_logic := '0';
    P31CTI	: in std_logic := '0';
    P31CTO	: out std_logic := '0';
    P31EI1	: in std_logic := '0';
    P31EI2	: in std_logic := '0';
    P31EI3	: in std_logic := '0';
    P31EI4	: in std_logic := '0';
    P31EI5	: in std_logic := '0';
    P31EI6	: in std_logic := '0';
    P31EI7	: in std_logic := '0';
    P31EI8	: in std_logic := '0';
    P31EL	: in std_logic := '0';
    P31ER	: in std_logic := '0';
    P31EO	: out std_logic := '0';
    P31RI	: in std_logic := '0';
    P31RL	: in std_logic := '0';
    P31RR	: in std_logic := '0';
    P31RO1	: out std_logic := '0';
    P31RO2	: out std_logic := '0';
    P31RO3	: out std_logic := '0';
    P31RO4	: out std_logic := '0';
    P31RO5	: out std_logic := '0';
    P31RO6	: out std_logic := '0';
    P31RO7	: out std_logic := '0';
    P31RO8	: out std_logic := '0';

    P32CI1	: in std_logic := '0';
    P32CL	: in std_logic := '0';
    P32CR	: in std_logic := '0';
    P32CO	: out std_logic := '0';
    P32CTI	: in std_logic := '0';
    P32CTO	: out std_logic := '0';
    P32EI1	: in std_logic := '0';
    P32EI2	: in std_logic := '0';
    P32EI3	: in std_logic := '0';
    P32EI4	: in std_logic := '0';
    P32EI5	: in std_logic := '0';
    P32EI6	: in std_logic := '0';
    P32EI7	: in std_logic := '0';
    P32EI8	: in std_logic := '0';
    P32EL	: in std_logic := '0';
    P32ER	: in std_logic := '0';
    P32EO	: out std_logic := '0';
    P32RI	: in std_logic := '0';
    P32RL	: in std_logic := '0';
    P32RR	: in std_logic := '0';
    P32RO1	: out std_logic := '0';
    P32RO2	: out std_logic := '0';
    P32RO3	: out std_logic := '0';
    P32RO4	: out std_logic := '0';
    P32RO5	: out std_logic := '0';
    P32RO6	: out std_logic := '0';
    P32RO7	: out std_logic := '0';
    P32RO8	: out std_logic := '0';

    P33CI1	: in std_logic := '0';
    P33CL	: in std_logic := '0';
    P33CR	: in std_logic := '0';
    P33CO	: out std_logic := '0';
    P33CTI	: in std_logic := '0';
    P33CTO	: out std_logic := '0';
    P33EI1	: in std_logic := '0';
    P33EI2	: in std_logic := '0';
    P33EI3	: in std_logic := '0';
    P33EI4	: in std_logic := '0';
    P33EI5	: in std_logic := '0';
    P33EI6	: in std_logic := '0';
    P33EI7	: in std_logic := '0';
    P33EI8	: in std_logic := '0';
    P33EL	: in std_logic := '0';
    P33ER	: in std_logic := '0';
    P33EO	: out std_logic := '0';
    P33RI	: in std_logic := '0';
    P33RL	: in std_logic := '0';
    P33RR	: in std_logic := '0';
    P33RO1	: out std_logic := '0';
    P33RO2	: out std_logic := '0';
    P33RO3	: out std_logic := '0';
    P33RO4	: out std_logic := '0';
    P33RO5	: out std_logic := '0';
    P33RO6	: out std_logic := '0';
    P33RO7	: out std_logic := '0';
    P33RO8	: out std_logic := '0';

    P34CI1	: in std_logic := '0';
    P34CL	: in std_logic := '0';
    P34CR	: in std_logic := '0';
    P34CO	: out std_logic := '0';
    P34CTI	: in std_logic := '0';
    P34CTO	: out std_logic := '0';
    P34EI1	: in std_logic := '0';
    P34EI2	: in std_logic := '0';
    P34EI3	: in std_logic := '0';
    P34EI4	: in std_logic := '0';
    P34EI5	: in std_logic := '0';
    P34EI6	: in std_logic := '0';
    P34EI7	: in std_logic := '0';
    P34EI8	: in std_logic := '0';
    P34EL	: in std_logic := '0';
    P34ER	: in std_logic := '0';
    P34EO	: out std_logic := '0';
    P34RI	: in std_logic := '0';
    P34RL	: in std_logic := '0';
    P34RR	: in std_logic := '0';
    P34RO1	: out std_logic := '0';
    P34RO2	: out std_logic := '0';
    P34RO3	: out std_logic := '0';
    P34RO4	: out std_logic := '0';
    P34RO5	: out std_logic := '0';
    P34RO6	: out std_logic := '0';
    P34RO7	: out std_logic := '0';
    P34RO8	: out std_logic := '0'
);
end component NX_IOM_U;

component NX_IOM_CONTROL_U is
generic (
    mode_side1        : integer := 0;
    div1         : bit_vector(2 downto 0) := "000";
    mode_side2        : integer := 0;
    div2         : bit_vector(2 downto 0) := "000";
    mode_side3        : integer := 0;
    div3         : bit_vector(2 downto 0) := "000";

    div_swrx1    : bit_vector(2 downto 0) := "000";
    div_swrx2    : bit_vector(2 downto 0) := "000";

    sel_ld_fck1  : bit_vector(1 downto 0) := "00";
    sel_ld_fck2  : bit_vector(1 downto 0) := "00";
    sel_ld_fck3  : bit_vector(1 downto 0) := "00";
    sel_sw_fck1  : bit_vector(1 downto 0) := "00";
    sel_sw_fck2  : bit_vector(1 downto 0) := "00";

    sel_dc_clk   : bit_vector(1 downto 0) := "00";

    inv_ld_sck1  : bit := '0';
    inv_ld_sck2  : bit := '0';
    inv_ld_sck3  : bit := '0';

    link_ld_12   : bit := '0';
    link_ld_23   : bit := '0';

    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';

    use_dc       : bit := '0';
    cal_delay1   : string := "";
    cal_delay2   : string := "";

    location     : string := ""
);
port (
    ALCK1	: in std_logic := '0';
    ALCK2	: in std_logic := '0';
    ALCK3	: in std_logic := '0';
    LDSCK1	: in std_logic := '0';
    LDSCK2	: in std_logic := '0';
    LDSCK3	: in std_logic := '0';
--  LDFCK1  : in    std_logic;	-- CONFIG
--  LDFCK2  : in    std_logic;	-- CONFIG
--  LDFCK3  : in    std_logic;	-- CONFIG
--  SWTX1CK : in    std_logic;	-- CONFIG
--  SWTX2CK : in    std_logic;	-- CONFIG
    SWRX1CK	: in std_logic := '0';
    SWRX2CK	: in std_logic := '0';
    FCK1	: in std_logic := '0';
    FCK2	: in std_logic := '0';
    FDCK	: in std_logic := '0';
    CCK	: in std_logic := '0';

    DQ1CI1	: in std_logic := '0';
    DQ1CI2	: in std_logic := '0';
    DQ1CI3	: in std_logic := '0';
    DQ1CI4	: in std_logic := '0';
    DQ1CI5	: in std_logic := '0';
    DQ1CI6	: in std_logic := '0';
    DQ1CI7	: in std_logic := '0';
    DQ1CI8	: in std_logic := '0';
    DQ2CI1	: in std_logic := '0';
    DQ2CI2	: in std_logic := '0';
    DQ2CI3	: in std_logic := '0';
    DQ2CI4	: in std_logic := '0';
    DQ2CI5	: in std_logic := '0';
    DQ2CI6	: in std_logic := '0';
    DQ2CI7	: in std_logic := '0';
    DQ2CI8	: in std_logic := '0';
    DQ3CI1	: in std_logic := '0';
    DQ3CI2	: in std_logic := '0';
    DQ3CI3	: in std_logic := '0';
    DQ3CI4	: in std_logic := '0';
    DQ3CI5	: in std_logic := '0';
    DQ3CI6	: in std_logic := '0';
    DQ3CI7	: in std_logic := '0';
    DQ3CI8	: in std_logic := '0';
    DQS1CI1	: in std_logic := '0';
    DQS1CI2	: in std_logic := '0';
    DQS1CI3	: in std_logic := '0';
    DQS1CI4	: in std_logic := '0';
    DQS1CI5	: in std_logic := '0';
    DQS1CI6	: in std_logic := '0';
    DQS1CI7	: in std_logic := '0';
    DQS1CI8	: in std_logic := '0';
    DQS2CI1	: in std_logic := '0';
    DQS2CI2	: in std_logic := '0';
    DQS2CI3	: in std_logic := '0';
    DQS2CI4	: in std_logic := '0';
    DQS2CI5	: in std_logic := '0';
    DQS2CI6	: in std_logic := '0';
    DQS2CI7	: in std_logic := '0';
    DQS2CI8	: in std_logic := '0';
    DQS3CI1	: in std_logic := '0';
    DQS3CI2	: in std_logic := '0';
    DQS3CI3	: in std_logic := '0';
    DQS3CI4	: in std_logic := '0';
    DQS3CI5	: in std_logic := '0';
    DQS3CI6	: in std_logic := '0';
    DQS3CI7	: in std_logic := '0';
    DQS3CI8	: in std_logic := '0';

    LD1RN	: in std_logic := '0';
    LD2RN	: in std_logic := '0';
    LD3RN	: in std_logic := '0';

    FA1	: in std_logic := '0';
    FA2	: in std_logic := '0';
    FA3	: in std_logic := '0';
    FA4	: in std_logic := '0';
    FA5	: in std_logic := '0';
    FA6	: in std_logic := '0';
    FZ	: in std_logic := '0';

    DCRN	: in std_logic := '0';
    LE	: in std_logic := '0';
    SE	: in std_logic := '0';

    DRI1	: in std_logic := '0';
    DRI2	: in std_logic := '0';
    DRI3	: in std_logic := '0';
    DRI4	: in std_logic := '0';
    DRI5	: in std_logic := '0';
    DRI6	: in std_logic := '0';
    DRA1	: in std_logic := '0';
    DRA2	: in std_logic := '0';
    DRA3	: in std_logic := '0';
    DRA4	: in std_logic := '0';

    DRO1CSN	: in std_logic := '0';
    DRO2CSN	: in std_logic := '0';
    DRO3CSN	: in std_logic := '0';
    DRI1CSN	: in std_logic := '0';
    DRI2CSN	: in std_logic := '0';
    DRI3CSN	: in std_logic := '0';
    DRDPA1CSN	: in std_logic := '0';
    DRDPA2CSN	: in std_logic := '0';
    DRDPA3CSN	: in std_logic := '0';
    DRCCSN	: in std_logic := '0';
    DRWDS	: in std_logic := '0';
    DRWEN	: in std_logic := '0';
    DRE	: in std_logic := '0';

    CA1P1	: in std_logic := '0';
    CA1P2	: in std_logic := '0';
    CA1P3	: in std_logic := '0';
    CA1P4	: in std_logic := '0';
    CA2P1	: in std_logic := '0';
    CA2P2	: in std_logic := '0';
    CA2P3	: in std_logic := '0';
    CA2P4	: in std_logic := '0';
    CA1N1	: in std_logic := '0';
    CA1N2	: in std_logic := '0';
    CA1N3	: in std_logic := '0';
    CA1N4	: in std_logic := '0';
    CA2N1	: in std_logic := '0';
    CA2N2	: in std_logic := '0';
    CA2N3	: in std_logic := '0';
    CA2N4	: in std_logic := '0';
    CA1T1	: in std_logic := '0';
    CA1T2	: in std_logic := '0';
    CA1T3	: in std_logic := '0';
    CA1T4	: in std_logic := '0';
    CA2T1	: in std_logic := '0';
    CA2T2	: in std_logic := '0';
    CA2T3	: in std_logic := '0';
    CA2T4	: in std_logic := '0';
    CA1D1	: in std_logic := '0';
    CA1D2	: in std_logic := '0';
    CA1D3	: in std_logic := '0';
    CA1D4	: in std_logic := '0';
    CA1D5	: in std_logic := '0';
    CA1D6	: in std_logic := '0';
    CA2D1	: in std_logic := '0';
    CA2D2	: in std_logic := '0';
    CA2D3	: in std_logic := '0';
    CA2D4	: in std_logic := '0';
    CA2D5	: in std_logic := '0';
    CA2D6	: in std_logic := '0';

    CKO1	: out std_logic := '0';
    CKO2	: out std_logic := '0';

    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0';
    AL1D	: out std_logic := '0';
    AL2D	: out std_logic := '0';
    AL3D	: out std_logic := '0';
    AL1T	: out std_logic := '0';
    AL2T	: out std_logic := '0';
    AL3T	: out std_logic := '0';
    DCL	: out std_logic := '0';
    DRO1	: out std_logic := '0';
    DRO2	: out std_logic := '0';
    DRO3	: out std_logic := '0';
    DRO4	: out std_logic := '0';
    DRO5	: out std_logic := '0';
    DRO6	: out std_logic := '0';

    LINK1	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK2	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK3	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK4	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK5	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK6	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK7	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK8	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK9	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK10	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK11	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK12	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK13	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK14	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK15	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK16	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK17	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK18	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK19	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK20	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK21	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK22	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK23	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK24	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK25	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK26	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK27	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK28	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK29	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK30	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK31	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK32	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK33	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0');
    LINK34	: inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0) := (others => '0')
);
end component NX_IOM_CONTROL_U;

component NX_PLL_L is
generic (
    location	      : string := "";
                      
    ref_intdiv        : integer   range 0 to 31 := 0;  -- 0 to 31  (%1 to %32)
    ref_osc_on        : bit := '0';                    -- 0: disabled - 1: enabled
                      
    cfg_use_pll       : std_logic:='1';                -- use or bypass PLL
                      
    ext_fbk_on        : bit := '0';                    -- 0: disabled - 1: enabled
                      
    fbk_intdiv        : integer   range 0 to 31 := 2;  -- 0 to 31  (%4 to %66 by step 2)
                      
    fbk_delay_on      : bit := '0';                    -- 0: no delay - 1: delay
    fbk_delay         : integer   range 0 to 63 := 0;  -- 0 to 63

    wfg_sync_pll_lock : bit := '0';                    -- 0: disabled - 1: enabled
    wfg_sync_cal_lock : bit := '0';                    -- 0: disabled - 1: enabled

    clk_outdivp1      : integer   range 0 to 7 := 0;   -- 0 to 7  P1 (2^n    : %1 to %128)
    clk_outdivp2      : integer   range 0 to 7 := 0;   -- 0 to 7  P2 (2^(n+1): %2 to %256)
    clk_outdivo1      : integer   range 0 to 7 := 0;   -- 0 to 7  O1 ((2n)+3 : %3 to  %17)
    clk_outdivp3o2    : integer   range 0 to 7 := 0    -- 0 to 7  P3 (2^(n+2): %4 to %512)
                                                       --         O2 ((2n)+5 : %5 to  %19)
);
port (
    REF	: in std_logic := '0';
    FBK	: in std_logic := '0';

    R	: in std_logic := '0';

    VCO	: out std_logic := '0';
    LDFO	: out std_logic := '0';
    REFO	: out std_logic := '0';

    DIVO1	: out std_logic := '0';
    DIVO2	: out std_logic := '0';

    DIVP1	: out std_logic := '0';
    DIVP2	: out std_logic := '0';
    DIVP3	: out std_logic := '0';
    OSC	: out std_logic := '0';

    PLL_LOCKED	: out std_logic := '0';
    CAL_LOCKED	: out std_logic := '0'
);
end component NX_PLL_L;

component NX_WFG_L is
generic (
    location    : string := "";
    wfg_edge    : bit := '0';                              -- 0: no invert / Rising
                                                           -- 1:    invert / Falling

    mode        : bit := '0';                              -- 0: no pattern - 1: pattern
    pattern_end : integer   range 0 to 15 := 1;            -- 0: to 15 (1 step to 16 steps)
    pattern     : bit_vector(0 to 15) := (others => '0');  -- pattern p0 ... p15

    delay_on    : bit := '0';                              -- 0: no delay - 1: delay
    delay       : integer   range 0 to 63 := 0             -- 0 to 63 (1 unit to 64 unit)
);
port (
    R	: in std_logic := '0';
    SI	: in std_logic := '0';
    ZI	: in std_logic := '0';
    RDY	: in std_logic := '1';
    SO	: out std_logic := '0';
    ZO	: out std_logic := '0'
);
end component NX_WFG_L;

component NX_PLL is
generic (
    location     : string := "";

    vco_range    : integer   range 0 to 2 := 0;   -- 0 to 3
    ref_div_on   : bit := '0';                    -- bypass :: %2
    fbk_div_on   : bit := '0';                    -- bypass :: %2
    ext_fbk_on   : bit := '0';                    -- 0: disabled - 1: enabled

    fbk_intdiv   : integer   range 1 to 31 := 2;  -- 0 to 31  (%1 to %32)

    fbk_delay_on : bit := '0';                    -- 0: no delay - 1: delay
    fbk_delay    : integer   range 0 to 63 := 0;  -- 0 to 63

    clk_outdiv1  : integer   range 0 to 7 := 0;   -- 0 to 7   (%1 to %2^7)
    clk_outdiv2  : integer   range 0 to 7 := 0;   -- 0 to 7   (%1 to %2^7)
    clk_outdiv3  : integer   range 0 to 7 := 0    -- 0 to 7   (%1 to %2^7)
);
port (
    REF	: in std_logic := '0';
    FBK	: in std_logic := '0';

    VCO	: out std_logic := '0';

    D1	: out std_logic := '0';
    D2	: out std_logic := '0';
    D3	: out std_logic := '0';
    OSC	: out std_logic := '0';

    RDY	: out std_logic := '0'
);
end component NX_PLL;

component NX_WFG is
generic (
    location    : string := "";

    wfg_edge    : bit := '0';                              -- 0: no invert / Rising
    mode        : bit := '0';                              -- 0: no pattern - 1: pattern

    pattern_end : integer   range 0 to 15 := 1;            -- 0: to 15 (1 step to 16 steps)
    pattern     : bit_vector(0 to 15) := (others => '0');  -- pattern p0 ... p15

    delay_on    : bit := '0';                              -- 0: no delay - 1: delay
    delay       : integer   range 0 to 63 := 0             -- 0 to 63 (1 unit to 64 unit)
);
port (
    SI	: in std_logic := '0';
    ZI	: in std_logic := '0';
    RDY	: in std_logic := '1';
    SO	: out std_logic := '0';
    ZO	: out std_logic := '0'
);
end component NX_WFG;

component NX_PLL_U is
generic (
        location     : string                 := "";               
        use_pll      : bit                    := '0';             -- Use the PLL
        pll_odf      : bit_vector(1 downto 0) := (others => '0'); -- Output division Factor
        pll_cpump    : bit_vector(3 downto 0) := (others => '0'); -- Set the charge pump factor
        pll_lpf_res  : bit_vector(3 downto 0) := (others => '0'); -- Set the resistances of the loop filter
        pll_lpf_cap  : bit_vector(3 downto 0) := (others => '0'); -- Set the capacitors of the loop filter
        pll_lock     : bit_vector(3 downto 0) := (others => '0'); -- Configuration of the frequency lock
        fbk_intdiv   : bit_vector(6 downto 0) := (others => '0'); -- Loop division Factor
        ref_intdiv   : bit_vector(4 downto 0) := (others => '0'); -- Reference Clock division Factor
        ref_osc_on   : bit                    := '0';             -- Reference Clock selection
        ext_fbk_on   : bit                    := '0';             -- Feedback Clock selection
        fbk_delay_on : bit                    := '0';             -- Add delay on the feedback clock
        fbk_delay    : bit_vector(5 downto 0) := (others => '0'); -- Delay on the feedback clock
        clk_outdiv1  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+3)
        clk_outdiv2  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+5)
        clk_outdiv3  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+7)
        clk_outdiv4  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+9)
        clk_outdivd1 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd2 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd3 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd4 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd5 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        use_cal      : bit                    := '0';             -- Use internal calibration
        clk_cal_sel  : bit_vector(1 downto 0) := "01";            -- Internal calibration clock selector
        cal_div      : bit_vector(3 downto 0) := "0111";          -- Division factor on Internal calibration clock
        cal_delay    : bit_vector(5 downto 0) := "011011"         -- Delay on internal calibration clock
    );
port (
    R	: in std_logic := '0';
    REF	: in std_logic := '0';
    FBK	: in std_logic := '0';
        -- Clock
    OSC	: out std_logic := '0';
    VCO	: out std_logic := '0';
    LDFO	: out std_logic := '0';
    REFO	: out std_logic := '0';
    CLK_DIV1	: out std_logic := '0';
    CLK_DIV2	: out std_logic := '0';
    CLK_DIV3	: out std_logic := '0';
    CLK_DIV4	: out std_logic := '0';
    CLK_DIVD1	: out std_logic := '0';
    CLK_DIVD2	: out std_logic := '0';
    CLK_DIVD3	: out std_logic := '0';
    CLK_DIVD4	: out std_logic := '0';
    CLK_DIVD5	: out std_logic := '0';
        -- Lock engine
    PLL_LOCKED	: out std_logic := '0';
    PLL_LOCKEDA	: out std_logic := '0';
        -- Calbration
    ARST_CAL	: in std_logic := '0';
    CLK_CAL	: in std_logic := '0';
    CLK_CAL_DIV	: out std_logic := '0';
    CAL_LOCKED	: out std_logic := '0';
    EXT_CAL_LOCKED	: in std_logic := '0';
    CAL1	: out std_logic := '0';
    CAL2	: out std_logic := '0';
    CAL3	: out std_logic := '0';
    CAL4	: out std_logic := '0';
    CAL5	: out std_logic := '0';
    EXT_CAL1	: in std_logic := '0';
    EXT_CAL2	: in std_logic := '0';
    EXT_CAL3	: in std_logic := '0';
    EXT_CAL4	: in std_logic := '0';
    EXT_CAL5	: in std_logic := '0'
    );
end component NX_PLL_U;

component NX_PLL_U_WRAP is
generic (
        location     : string                 := ""; 
        use_pll      : bit                    := '0';             -- Use the PLL
        pll_odf      : bit_vector(1 downto 0) := (others => '0'); -- Output division Factor
        pll_cpump    : bit_vector(3 downto 0) := (others => '0'); -- Set the charge pump factor
        pll_lpf_res  : bit_vector(3 downto 0) := (others => '0'); -- Set the resistances of the loop filter
        pll_lpf_cap  : bit_vector(3 downto 0) := (others => '0'); -- Set the capacitors of the loop filter
        pll_lock     : bit_vector(3 downto 0) := (others => '0'); -- Configuration of the frequency lock
        fbk_intdiv   : bit_vector(6 downto 0) := (others => '0'); -- Loop division Factor
        ref_intdiv   : bit_vector(4 downto 0) := (others => '0'); -- Reference Clock division Factor
        ref_osc_on   : bit                    := '0';             -- Reference Clock selection
        ext_fbk_on   : bit                    := '0';             -- Feedback Clock selection
        fbk_delay_on : bit                    := '0';             -- Add delay on the feedback clock
        fbk_delay    : bit_vector(5 downto 0) := (others => '0'); -- Delay on the feedback clock
        clk_outdiv1  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+3)
        clk_outdiv2  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+5)
        clk_outdiv3  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+7)
        clk_outdiv4  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+9)
        clk_outdivd1 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd2 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd3 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd4 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd5 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        use_cal      : bit                    := '0';             -- Use internal calibration
        clk_cal_sel  : bit_vector(1 downto 0) := "01";            -- Internal calibration clock selector
        cal_div      : bit_vector(3 downto 0) := "0111";          -- Division factor on Internal calibration clock
        cal_delay    : bit_vector(5 downto 0) := "011011"         -- Delay on internal calibration clock
    );
port (
    R	: in std_logic := '0';
    REF	: in std_logic := '0';
    FBK	: in std_logic := '0';
        -- Clock
    OSC	: out std_logic := '0';
    VCO	: out std_logic := '0';
    LDFO	: out std_logic := '0';
    REFO	: out std_logic := '0';
    CLK_DIV	: out std_logic_vector(3 downto 0); -- 0 : 1/(N+3); 1 : 1/(N+5); 2 : 1/(N+7) := (others => '0');
    CLK_DIVD	: out std_logic_vector(4 downto 0) := (others => '0');
        -- Lock engine
    PLL_LOCKED	: out std_logic := '0';
    PLL_LOCKEDA	: out std_logic := '0';
        -- Calibration
    ARST_CAL	: in std_logic := '0';
    CLK_CAL	: in std_logic := '0';
    CLK_CAL_DIV	: out std_logic := '0';
    CAL_LOCKED	: out std_logic := '0';
    EXT_CAL_LOCKED	: in std_logic := '0';
    CAL	: out std_logic_vector(4 downto 0) := (others => '0');
    EXT_CAL	: in std_logic_vector(4 downto 0) := (others => '0')
    );
end component NX_PLL_U_WRAP;

component NX_WFG_U is
generic (
        location             : string := "";
        wfg_edge             : bit                   := '0'; -- 0: no invert / Rising
        reset_on_pll_lock_n  : bit                   := '0';
        reset_on_pll_locka_n : bit                   := '0';
        reset_on_cal_lock_n  : bit                   := '0';

        mode                 : integer range 0 to 2 := 0;                                   -- 0: no pattern - 1: pattern - 2: diviseur
        pattern              : bit_vector(0 to 15)   := b"0000000000000000"; -- pattern p0 ... p15
        pattern_end          : integer range 0 to 15 := 0;                   -- max pattern length. Set to 0 to use divider/bypass instead of pattern
        div_ratio            : integer range 0 to 2047 := 0;                   -- divisor ratio
        delay_on             : bit                   := '0';                 -- 0: no delay - 1: delay
        delay                : integer range 0 to 63 := 0                    -- 0 to 63 (1 unit to 32 unit)
    );
port (
    R	: in std_logic := '0';
    SI	: in std_logic := '0';
    ZI	: in std_logic := '0';
    SO	: out std_logic := '0';
    ZO	: out std_logic := '0'
    );
end component NX_WFG_U;

component NX_R5_L is
port (
    -- Inputs
    A_CKEM_I	: in std_logic := '0';
    A_CKEP_I	: in std_logic := '0';
    A_CKES_I	: in std_logic := '0';

    AR_A_I32	: in std_logic := '0';
    AR_A_I31	: in std_logic := '0';
    AR_A_I30	: in std_logic := '0';
    AR_A_I29	: in std_logic := '0';
    AR_A_I28	: in std_logic := '0';
    AR_A_I27	: in std_logic := '0';
    AR_A_I26	: in std_logic := '0';
    AR_A_I25	: in std_logic := '0';
    AR_A_I24	: in std_logic := '0';
    AR_A_I23	: in std_logic := '0';
    AR_A_I22	: in std_logic := '0';
    AR_A_I21	: in std_logic := '0';
    AR_A_I20	: in std_logic := '0';
    AR_A_I19	: in std_logic := '0';
    AR_A_I18	: in std_logic := '0';
    AR_A_I17	: in std_logic := '0';
    AR_A_I16	: in std_logic := '0';
    AR_A_I15	: in std_logic := '0';
    AR_A_I14	: in std_logic := '0';
    AR_A_I13	: in std_logic := '0';
    AR_A_I12	: in std_logic := '0';
    AR_A_I11	: in std_logic := '0';
    AR_A_I10	: in std_logic := '0';
    AR_A_I9	: in std_logic := '0';
    AR_A_I8	: in std_logic := '0';
    AR_A_I7	: in std_logic := '0';
    AR_A_I6	: in std_logic := '0';
    AR_A_I5	: in std_logic := '0';
    AR_A_I4	: in std_logic := '0';
    AR_A_I3	: in std_logic := '0';
    AR_A_I2	: in std_logic := '0';
    AR_A_I1	: in std_logic := '0';

    AR_BU_I2	: in std_logic := '0';
    AR_BU_I1	: in std_logic := '0';

    AR_CH_I4	: in std_logic := '0';
    AR_CH_I3	: in std_logic := '0';
    AR_CH_I2	: in std_logic := '0';
    AR_CH_I1	: in std_logic := '0';

    AR_IDS_I8	: in std_logic := '0';
    AR_IDS_I7	: in std_logic := '0';
    AR_IDS_I6	: in std_logic := '0';
    AR_IDS_I5	: in std_logic := '0';
    AR_IDS_I4	: in std_logic := '0';
    AR_IDS_I3	: in std_logic := '0';
    AR_IDS_I2	: in std_logic := '0';
    AR_IDS_I1	: in std_logic := '0';

    AR_LE_I4	: in std_logic := '0';
    AR_LE_I3	: in std_logic := '0';
    AR_LE_I2	: in std_logic := '0';
    AR_LE_I1	: in std_logic := '0';

    AR_LK_I2	: in std_logic := '0';
    AR_LK_I1	: in std_logic := '0';

    AR_PR_I3	: in std_logic := '0';
    AR_PR_I2	: in std_logic := '0';
    AR_PR_I1	: in std_logic := '0';

    AR_RYM_I	: in std_logic := '0';
    AR_RYP_I	: in std_logic := '0';

    AR_SZ_I3	: in std_logic := '0';
    AR_SZ_I2	: in std_logic := '0';
    AR_SZ_I1	: in std_logic := '0';

    AR_VD_I	: in std_logic := '0';
    AT_RS_I	: in std_logic := '0';

    AW_A_I32	: in std_logic := '0';
    AW_A_I31	: in std_logic := '0';
    AW_A_I30	: in std_logic := '0';
    AW_A_I29	: in std_logic := '0';
    AW_A_I28	: in std_logic := '0';
    AW_A_I27	: in std_logic := '0';
    AW_A_I26	: in std_logic := '0';
    AW_A_I25	: in std_logic := '0';
    AW_A_I24	: in std_logic := '0';
    AW_A_I23	: in std_logic := '0';
    AW_A_I22	: in std_logic := '0';
    AW_A_I21	: in std_logic := '0';
    AW_A_I20	: in std_logic := '0';
    AW_A_I19	: in std_logic := '0';
    AW_A_I18	: in std_logic := '0';
    AW_A_I17	: in std_logic := '0';
    AW_A_I16	: in std_logic := '0';
    AW_A_I15	: in std_logic := '0';
    AW_A_I14	: in std_logic := '0';
    AW_A_I13	: in std_logic := '0';
    AW_A_I12	: in std_logic := '0';
    AW_A_I11	: in std_logic := '0';
    AW_A_I10	: in std_logic := '0';
    AW_A_I9	: in std_logic := '0';
    AW_A_I8	: in std_logic := '0';
    AW_A_I7	: in std_logic := '0';
    AW_A_I6	: in std_logic := '0';
    AW_A_I5	: in std_logic := '0';
    AW_A_I4	: in std_logic := '0';
    AW_A_I3	: in std_logic := '0';
    AW_A_I2	: in std_logic := '0';
    AW_A_I1	: in std_logic := '0';

    AW_BU_I2	: in std_logic := '0';
    AW_BU_I1	: in std_logic := '0';

    AW_CH_I4	: in std_logic := '0';
    AW_CH_I3	: in std_logic := '0';
    AW_CH_I2	: in std_logic := '0';
    AW_CH_I1	: in std_logic := '0';

    AW_IDS_I8	: in std_logic := '0';
    AW_IDS_I7	: in std_logic := '0';
    AW_IDS_I6	: in std_logic := '0';
    AW_IDS_I5	: in std_logic := '0';
    AW_IDS_I4	: in std_logic := '0';
    AW_IDS_I3	: in std_logic := '0';
    AW_IDS_I2	: in std_logic := '0';
    AW_IDS_I1	: in std_logic := '0';

    AW_LE_I4	: in std_logic := '0';
    AW_LE_I3	: in std_logic := '0';
    AW_LE_I2	: in std_logic := '0';
    AW_LE_I1	: in std_logic := '0';

    AW_LK_I2	: in std_logic := '0';
    AW_LK_I1	: in std_logic := '0';

    AW_PR_I3	: in std_logic := '0';
    AW_PR_I2	: in std_logic := '0';
    AW_PR_I1	: in std_logic := '0';

    AW_RYM_I	: in std_logic := '0';
    AW_RYP_I	: in std_logic := '0';

    AW_SZ_I3	: in std_logic := '0';
    AW_SZ_I2	: in std_logic := '0';
    AW_SZ_I1	: in std_logic := '0';

    AW_VD_I	: in std_logic := '0';

    B_IDM_I4	: in std_logic := '0';
    B_IDM_I3	: in std_logic := '0';
    B_IDM_I2	: in std_logic := '0';
    B_IDM_I1	: in std_logic := '0';

    B_IDP_I4	: in std_logic := '0';
    B_IDP_I3	: in std_logic := '0';
    B_IDP_I2	: in std_logic := '0';
    B_IDP_I1	: in std_logic := '0';

    B_RDY_I	: in std_logic := '0';

    B_RSPM_I2	: in std_logic := '0';
    B_RSPM_I1	: in std_logic := '0';

    B_RSPP_I2	: in std_logic := '0';
    B_RSPP_I1	: in std_logic := '0';

    B_VDM_I	: in std_logic := '0';
    B_VDP_I	: in std_logic := '0';

--    CAL_I5        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I4        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I3        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I2        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I1        : in  std_logic; --  calibration   5   [0:4]

    CDB_PW_I	: in std_logic := '0';
    CDB_RS_I	: in std_logic := '0';
    CFG_EE_I	: in std_logic := '0';
    CFG_IE_I	: in std_logic := '0';
    CFG_NM_I	: in std_logic := '0';
    CK_I	: in std_logic := '0';
--    CK_DR_I       : in  std_logic; --  clock_dr      1
    CS_PW_I	: in std_logic := '0';
    DB_E_I	: in std_logic := '0';
    DB_NCK_I	: in std_logic := '0';

    DB_RA_I20	: in std_logic := '0';
    DB_RA_I19	: in std_logic := '0';
    DB_RA_I18	: in std_logic := '0';
    DB_RA_I17	: in std_logic := '0';
    DB_RA_I16	: in std_logic := '0';
    DB_RA_I15	: in std_logic := '0';
    DB_RA_I14	: in std_logic := '0';
    DB_RA_I13	: in std_logic := '0';
    DB_RA_I12	: in std_logic := '0';
    DB_RA_I11	: in std_logic := '0';
    DB_RA_I10	: in std_logic := '0';
    DB_RA_I9	: in std_logic := '0';
    DB_RA_I8	: in std_logic := '0';
    DB_RA_I7	: in std_logic := '0';
    DB_RA_I6	: in std_logic := '0';
    DB_RA_I5	: in std_logic := '0';
    DB_RA_I4	: in std_logic := '0';
    DB_RA_I3	: in std_logic := '0';
    DB_RA_I2	: in std_logic := '0';
    DB_RA_I1	: in std_logic := '0';

    DB_RAV_I	: in std_logic := '0';

    DB_SA_I20	: in std_logic := '0';
    DB_SA_I19	: in std_logic := '0';
    DB_SA_I18	: in std_logic := '0';
    DB_SA_I17	: in std_logic := '0';
    DB_SA_I16	: in std_logic := '0';
    DB_SA_I15	: in std_logic := '0';
    DB_SA_I14	: in std_logic := '0';
    DB_SA_I13	: in std_logic := '0';
    DB_SA_I12	: in std_logic := '0';
    DB_SA_I11	: in std_logic := '0';
    DB_SA_I10	: in std_logic := '0';
    DB_SA_I9	: in std_logic := '0';
    DB_SA_I8	: in std_logic := '0';
    DB_SA_I7	: in std_logic := '0';
    DB_SA_I6	: in std_logic := '0';
    DB_SA_I5	: in std_logic := '0';
    DB_SA_I4	: in std_logic := '0';
    DB_SA_I3	: in std_logic := '0';
    DB_SA_I2	: in std_logic := '0';
    DB_SA_I1	: in std_logic := '0';

    DB_SAV_I	: in std_logic := '0';
    DEV_E_I	: in std_logic := '0';

    DFTS_I8	: in std_logic := '0';
    DFTS_I7	: in std_logic := '0';
    DFTS_I6	: in std_logic := '0';
    DFTS_I5	: in std_logic := '0';
    DFTS_I4	: in std_logic := '0';
    DFTS_I3	: in std_logic := '0';
    DFTS_I2	: in std_logic := '0';
    DFTS_I1	: in std_logic := '0';

    E_DB_I	: in std_logic := '0';
    ERR_R_I	: in std_logic := '0';
    EVENT_I	: in std_logic := '0';

    GID_I4	: in std_logic := '0';
    GID_I3	: in std_logic := '0';
    GID_I2	: in std_logic := '0';
    GID_I1	: in std_logic := '0';

    INIT_P_I	: in std_logic := '0';
    INIT_R_I	: in std_logic := '0';
    LOC_R_I	: in std_logic := '0';
--    LBK_E_I       : in  std_logic; --  loopback_en   1
--    LBK_MX_I      : in  std_logic; --  loopback_mux  1

--    MODE1_I3      : in  std_logic; --  mode1         3   [0:2]
--    MODE1_I2      : in  std_logic; --  mode1         3   [0:2]
--    MODE1_I1      : in  std_logic; --  mode1         3   [0:2]

--    MODE2_I3      : in  std_logic; --  mode2         3   [0:2]
--    MODE2_I2      : in  std_logic; --  mode2         3   [0:2]
--    MODE2_I1      : in  std_logic; --  mode2         3   [0:2]

--    MODE3_I3      : in  std_logic; --  mode3         3   [0:2]
--    MODE3_I2      : in  std_logic; --  mode3         3   [0:2]
--    MODE3_I1      : in  std_logic; --  mode3         3   [0:2]

    NCPUH_I	: in std_logic := '0';
    NET_RS_I	: in std_logic := '0';
    N_FIQ_I	: in std_logic := '0';
    N_IDE_I	: in std_logic := '0';
    N_IRQ_I	: in std_logic := '0';
    N_PRS_I	: in std_logic := '0';
    N_RS_I	: in std_logic := '0';
    N_SPRS_I	: in std_logic := '0';
    N_TRS_I	: in std_logic := '0';

    P_A_I29	: in std_logic := '0';
    P_A_I28	: in std_logic := '0';
    P_A_I27	: in std_logic := '0';
    P_A_I26	: in std_logic := '0';
    P_A_I25	: in std_logic := '0';
    P_A_I24	: in std_logic := '0';
    P_A_I23	: in std_logic := '0';
    P_A_I22	: in std_logic := '0';
    P_A_I21	: in std_logic := '0';
    P_A_I20	: in std_logic := '0';
    P_A_I19	: in std_logic := '0';
    P_A_I18	: in std_logic := '0';
    P_A_I17	: in std_logic := '0';
    P_A_I16	: in std_logic := '0';
    P_A_I15	: in std_logic := '0';
    P_A_I14	: in std_logic := '0';
    P_A_I13	: in std_logic := '0';
    P_A_I12	: in std_logic := '0';
    P_A_I11	: in std_logic := '0';
    P_A_I10	: in std_logic := '0';
    P_A_I9	: in std_logic := '0';
    P_A_I8	: in std_logic := '0';
    P_A_I7	: in std_logic := '0';
    P_A_I6	: in std_logic := '0';
    P_A_I5	: in std_logic := '0';
    P_A_I4	: in std_logic := '0';
    P_A_I3	: in std_logic := '0';
    P_A_I2	: in std_logic := '0';
    P_A_I1	: in std_logic := '0';

    P_ECC_I	: in std_logic := '0';
    PLVL_I	: in std_logic := '0';
    P_CK_E_I	: in std_logic := '0';
    P_CK_I	: in std_logic := '0';
    P_E_I	: in std_logic := '0';

    PPV_BS_I20	: in std_logic := '0';
    PPV_BS_I19	: in std_logic := '0';
    PPV_BS_I18	: in std_logic := '0';
    PPV_BS_I17	: in std_logic := '0';
    PPV_BS_I16	: in std_logic := '0';
    PPV_BS_I15	: in std_logic := '0';
    PPV_BS_I14	: in std_logic := '0';
    PPV_BS_I13	: in std_logic := '0';
    PPV_BS_I12	: in std_logic := '0';
    PPV_BS_I11	: in std_logic := '0';
    PPV_BS_I10	: in std_logic := '0';
    PPV_BS_I9	: in std_logic := '0';
    PPV_BS_I8	: in std_logic := '0';
    PPV_BS_I7	: in std_logic := '0';
    PPV_BS_I6	: in std_logic := '0';
    PPV_BS_I5	: in std_logic := '0';
    PPV_BS_I4	: in std_logic := '0';
    PPV_BS_I3	: in std_logic := '0';
    PPV_BS_I2	: in std_logic := '0';
    PPV_BS_I1	: in std_logic := '0';

    PPV_SZ_I5	: in std_logic := '0';
    PPV_SZ_I4	: in std_logic := '0';
    PPV_SZ_I3	: in std_logic := '0';
    PPV_SZ_I2	: in std_logic := '0';
    PPV_SZ_I1	: in std_logic := '0';

    PPX_BS_I20	: in std_logic := '0';
    PPX_BS_I19	: in std_logic := '0';
    PPX_BS_I18	: in std_logic := '0';
    PPX_BS_I17	: in std_logic := '0';
    PPX_BS_I16	: in std_logic := '0';
    PPX_BS_I15	: in std_logic := '0';
    PPX_BS_I14	: in std_logic := '0';
    PPX_BS_I13	: in std_logic := '0';
    PPX_BS_I12	: in std_logic := '0';
    PPX_BS_I11	: in std_logic := '0';
    PPX_BS_I10	: in std_logic := '0';
    PPX_BS_I9	: in std_logic := '0';
    PPX_BS_I8	: in std_logic := '0';
    PPX_BS_I7	: in std_logic := '0';
    PPX_BS_I6	: in std_logic := '0';
    PPX_BS_I5	: in std_logic := '0';
    PPX_BS_I4	: in std_logic := '0';
    PPX_BS_I3	: in std_logic := '0';
    PPX_BS_I2	: in std_logic := '0';
    PPX_BS_I1	: in std_logic := '0';

    PPX_SZ_I5	: in std_logic := '0';
    PPX_SZ_I4	: in std_logic := '0';
    PPX_SZ_I3	: in std_logic := '0';
    PPX_SZ_I2	: in std_logic := '0';
    PPX_SZ_I1	: in std_logic := '0';

    P_RS_I	: in std_logic := '0';
    P_SEL_I	: in std_logic := '0';

    PW_D_I32	: in std_logic := '0';
    PW_D_I31	: in std_logic := '0';
    PW_D_I30	: in std_logic := '0';
    PW_D_I29	: in std_logic := '0';
    PW_D_I28	: in std_logic := '0';
    PW_D_I27	: in std_logic := '0';
    PW_D_I26	: in std_logic := '0';
    PW_D_I25	: in std_logic := '0';
    PW_D_I24	: in std_logic := '0';
    PW_D_I23	: in std_logic := '0';
    PW_D_I22	: in std_logic := '0';
    PW_D_I21	: in std_logic := '0';
    PW_D_I20	: in std_logic := '0';
    PW_D_I19	: in std_logic := '0';
    PW_D_I18	: in std_logic := '0';
    PW_D_I17	: in std_logic := '0';
    PW_D_I16	: in std_logic := '0';
    PW_D_I15	: in std_logic := '0';
    PW_D_I14	: in std_logic := '0';
    PW_D_I13	: in std_logic := '0';
    PW_D_I12	: in std_logic := '0';
    PW_D_I11	: in std_logic := '0';
    PW_D_I10	: in std_logic := '0';
    PW_D_I9	: in std_logic := '0';
    PW_D_I8	: in std_logic := '0';
    PW_D_I7	: in std_logic := '0';
    PW_D_I6	: in std_logic := '0';
    PW_D_I5	: in std_logic := '0';
    PW_D_I4	: in std_logic := '0';
    PW_D_I3	: in std_logic := '0';
    PW_D_I2	: in std_logic := '0';
    PW_D_I1	: in std_logic := '0';

    PW_I	: in std_logic := '0';

    RAMCTL_I8	: in std_logic := '0';
    RAMCTL_I7	: in std_logic := '0';
    RAMCTL_I6	: in std_logic := '0';
    RAMCTL_I5	: in std_logic := '0';
    RAMCTL_I4	: in std_logic := '0';
    RAMCTL_I3	: in std_logic := '0';
    RAMCTL_I2	: in std_logic := '0';
    RAMCTL_I1	: in std_logic := '0';

    R_DM_I64	: in std_logic := '0';
    R_DM_I63	: in std_logic := '0';
    R_DM_I62	: in std_logic := '0';
    R_DM_I61	: in std_logic := '0';
    R_DM_I60	: in std_logic := '0';
    R_DM_I59	: in std_logic := '0';
    R_DM_I58	: in std_logic := '0';
    R_DM_I57	: in std_logic := '0';
    R_DM_I56	: in std_logic := '0';
    R_DM_I55	: in std_logic := '0';
    R_DM_I54	: in std_logic := '0';
    R_DM_I53	: in std_logic := '0';
    R_DM_I52	: in std_logic := '0';
    R_DM_I51	: in std_logic := '0';
    R_DM_I50	: in std_logic := '0';
    R_DM_I49	: in std_logic := '0';
    R_DM_I48	: in std_logic := '0';
    R_DM_I47	: in std_logic := '0';
    R_DM_I46	: in std_logic := '0';
    R_DM_I45	: in std_logic := '0';
    R_DM_I44	: in std_logic := '0';
    R_DM_I43	: in std_logic := '0';
    R_DM_I42	: in std_logic := '0';
    R_DM_I41	: in std_logic := '0';
    R_DM_I40	: in std_logic := '0';
    R_DM_I39	: in std_logic := '0';
    R_DM_I38	: in std_logic := '0';
    R_DM_I37	: in std_logic := '0';
    R_DM_I36	: in std_logic := '0';
    R_DM_I35	: in std_logic := '0';
    R_DM_I34	: in std_logic := '0';
    R_DM_I33	: in std_logic := '0';
    R_DM_I32	: in std_logic := '0';
    R_DM_I31	: in std_logic := '0';
    R_DM_I30	: in std_logic := '0';
    R_DM_I29	: in std_logic := '0';
    R_DM_I28	: in std_logic := '0';
    R_DM_I27	: in std_logic := '0';
    R_DM_I26	: in std_logic := '0';
    R_DM_I25	: in std_logic := '0';
    R_DM_I24	: in std_logic := '0';
    R_DM_I23	: in std_logic := '0';
    R_DM_I22	: in std_logic := '0';
    R_DM_I21	: in std_logic := '0';
    R_DM_I20	: in std_logic := '0';
    R_DM_I19	: in std_logic := '0';
    R_DM_I18	: in std_logic := '0';
    R_DM_I17	: in std_logic := '0';
    R_DM_I16	: in std_logic := '0';
    R_DM_I15	: in std_logic := '0';
    R_DM_I14	: in std_logic := '0';
    R_DM_I13	: in std_logic := '0';
    R_DM_I12	: in std_logic := '0';
    R_DM_I11	: in std_logic := '0';
    R_DM_I10	: in std_logic := '0';
    R_DM_I9	: in std_logic := '0';
    R_DM_I8	: in std_logic := '0';
    R_DM_I7	: in std_logic := '0';
    R_DM_I6	: in std_logic := '0';
    R_DM_I5	: in std_logic := '0';
    R_DM_I4	: in std_logic := '0';
    R_DM_I3	: in std_logic := '0';
    R_DM_I2	: in std_logic := '0';
    R_DM_I1	: in std_logic := '0';

    R_DP_I32	: in std_logic := '0';
    R_DP_I31	: in std_logic := '0';
    R_DP_I30	: in std_logic := '0';
    R_DP_I29	: in std_logic := '0';
    R_DP_I28	: in std_logic := '0';
    R_DP_I27	: in std_logic := '0';
    R_DP_I26	: in std_logic := '0';
    R_DP_I25	: in std_logic := '0';
    R_DP_I24	: in std_logic := '0';
    R_DP_I23	: in std_logic := '0';
    R_DP_I22	: in std_logic := '0';
    R_DP_I21	: in std_logic := '0';
    R_DP_I20	: in std_logic := '0';
    R_DP_I19	: in std_logic := '0';
    R_DP_I18	: in std_logic := '0';
    R_DP_I17	: in std_logic := '0';
    R_DP_I16	: in std_logic := '0';
    R_DP_I15	: in std_logic := '0';
    R_DP_I14	: in std_logic := '0';
    R_DP_I13	: in std_logic := '0';
    R_DP_I12	: in std_logic := '0';
    R_DP_I11	: in std_logic := '0';
    R_DP_I10	: in std_logic := '0';
    R_DP_I9	: in std_logic := '0';
    R_DP_I8	: in std_logic := '0';
    R_DP_I7	: in std_logic := '0';
    R_DP_I6	: in std_logic := '0';
    R_DP_I5	: in std_logic := '0';
    R_DP_I4	: in std_logic := '0';
    R_DP_I3	: in std_logic := '0';
    R_DP_I2	: in std_logic := '0';
    R_DP_I1	: in std_logic := '0';

--    RDY_I3        : in  std_logic; --  ready         3   [0:2]
--    RDY_I2        : in  std_logic; --  ready         3   [0:2]
--    RDY_I1        : in  std_logic; --  ready         3   [0:2]

    R_IDM_I4	: in std_logic := '0';
    R_IDM_I3	: in std_logic := '0';
    R_IDM_I2	: in std_logic := '0';
    R_IDM_I1	: in std_logic := '0';

    R_IDP_I4	: in std_logic := '0';
    R_IDP_I3	: in std_logic := '0';
    R_IDP_I2	: in std_logic := '0';
    R_IDP_I1	: in std_logic := '0';

    R_LSTM_I	: in std_logic := '0';
    R_LSTP_I	: in std_logic := '0';
    R_RDY_I	: in std_logic := '0';

    R_RSPM_I2	: in std_logic := '0';
    R_RSPM_I1	: in std_logic := '0';

    R_RSPP_I2	: in std_logic := '0';
    R_RSPP_I1	: in std_logic := '0';

    RS_BYP_I	: in std_logic := '0';
    R_VDM_I	: in std_logic := '0';
    R_VDP_I	: in std_logic := '0';
--    SCAN_E_I      : in  std_logic; --  scan_en       1
    SE_I	: in std_logic := '0';
--    SHF_DR_I      : in  std_logic; --  shift_dr      1
--    SH_I          : in  std_logic; --  shin          1
    SW_CK_I	: in std_logic := '0';
    SW_DI_I	: in std_logic := '0';
    T_DI_I	: in std_logic := '0';
    TE_INI_I	: in std_logic := '0';
--    TEST_E_I      : in  std_logic; --  test_en       1
--    UPD_DR_I      : in  std_logic; --  update_dr     1
    VINI_I	: in std_logic := '0';

    W_D_I64	: in std_logic := '0';
    W_D_I63	: in std_logic := '0';
    W_D_I62	: in std_logic := '0';
    W_D_I61	: in std_logic := '0';
    W_D_I60	: in std_logic := '0';
    W_D_I59	: in std_logic := '0';
    W_D_I58	: in std_logic := '0';
    W_D_I57	: in std_logic := '0';
    W_D_I56	: in std_logic := '0';
    W_D_I55	: in std_logic := '0';
    W_D_I54	: in std_logic := '0';
    W_D_I53	: in std_logic := '0';
    W_D_I52	: in std_logic := '0';
    W_D_I51	: in std_logic := '0';
    W_D_I50	: in std_logic := '0';
    W_D_I49	: in std_logic := '0';
    W_D_I48	: in std_logic := '0';
    W_D_I47	: in std_logic := '0';
    W_D_I46	: in std_logic := '0';
    W_D_I45	: in std_logic := '0';
    W_D_I44	: in std_logic := '0';
    W_D_I43	: in std_logic := '0';
    W_D_I42	: in std_logic := '0';
    W_D_I41	: in std_logic := '0';
    W_D_I40	: in std_logic := '0';
    W_D_I39	: in std_logic := '0';
    W_D_I38	: in std_logic := '0';
    W_D_I37	: in std_logic := '0';
    W_D_I36	: in std_logic := '0';
    W_D_I35	: in std_logic := '0';
    W_D_I34	: in std_logic := '0';
    W_D_I33	: in std_logic := '0';
    W_D_I32	: in std_logic := '0';
    W_D_I31	: in std_logic := '0';
    W_D_I30	: in std_logic := '0';
    W_D_I29	: in std_logic := '0';
    W_D_I28	: in std_logic := '0';
    W_D_I27	: in std_logic := '0';
    W_D_I26	: in std_logic := '0';
    W_D_I25	: in std_logic := '0';
    W_D_I24	: in std_logic := '0';
    W_D_I23	: in std_logic := '0';
    W_D_I22	: in std_logic := '0';
    W_D_I21	: in std_logic := '0';
    W_D_I20	: in std_logic := '0';
    W_D_I19	: in std_logic := '0';
    W_D_I18	: in std_logic := '0';
    W_D_I17	: in std_logic := '0';
    W_D_I16	: in std_logic := '0';
    W_D_I15	: in std_logic := '0';
    W_D_I14	: in std_logic := '0';
    W_D_I13	: in std_logic := '0';
    W_D_I12	: in std_logic := '0';
    W_D_I11	: in std_logic := '0';
    W_D_I10	: in std_logic := '0';
    W_D_I9	: in std_logic := '0';
    W_D_I8	: in std_logic := '0';
    W_D_I7	: in std_logic := '0';
    W_D_I6	: in std_logic := '0';
    W_D_I5	: in std_logic := '0';
    W_D_I4	: in std_logic := '0';
    W_D_I3	: in std_logic := '0';
    W_D_I2	: in std_logic := '0';
    W_D_I1	: in std_logic := '0';

    W_IDS_I8	: in std_logic := '0';
    W_IDS_I7	: in std_logic := '0';
    W_IDS_I6	: in std_logic := '0';
    W_IDS_I5	: in std_logic := '0';
    W_IDS_I4	: in std_logic := '0';
    W_IDS_I3	: in std_logic := '0';
    W_IDS_I2	: in std_logic := '0';
    W_IDS_I1	: in std_logic := '0';

    W_LST_I	: in std_logic := '0';
    W_RYM_I	: in std_logic := '0';
    W_RYP_I	: in std_logic := '0';

    W_SBS_I8	: in std_logic := '0';
    W_SBS_I7	: in std_logic := '0';
    W_SBS_I6	: in std_logic := '0';
    W_SBS_I5	: in std_logic := '0';
    W_SBS_I4	: in std_logic := '0';
    W_SBS_I3	: in std_logic := '0';
    W_SBS_I2	: in std_logic := '0';
    W_SBS_I1	: in std_logic := '0';

    W_VD_I	: in std_logic := '0';

    -- Outputs
    AR_AM_O32	: out std_logic := '0';
    AR_AM_O31	: out std_logic := '0';
    AR_AM_O30	: out std_logic := '0';
    AR_AM_O29	: out std_logic := '0';
    AR_AM_O28	: out std_logic := '0';
    AR_AM_O27	: out std_logic := '0';
    AR_AM_O26	: out std_logic := '0';
    AR_AM_O25	: out std_logic := '0';
    AR_AM_O24	: out std_logic := '0';
    AR_AM_O23	: out std_logic := '0';
    AR_AM_O22	: out std_logic := '0';
    AR_AM_O21	: out std_logic := '0';
    AR_AM_O20	: out std_logic := '0';
    AR_AM_O19	: out std_logic := '0';
    AR_AM_O18	: out std_logic := '0';
    AR_AM_O17	: out std_logic := '0';
    AR_AM_O16	: out std_logic := '0';
    AR_AM_O15	: out std_logic := '0';
    AR_AM_O14	: out std_logic := '0';
    AR_AM_O13	: out std_logic := '0';
    AR_AM_O12	: out std_logic := '0';
    AR_AM_O11	: out std_logic := '0';
    AR_AM_O10	: out std_logic := '0';
    AR_AM_O9	: out std_logic := '0';
    AR_AM_O8	: out std_logic := '0';
    AR_AM_O7	: out std_logic := '0';
    AR_AM_O6	: out std_logic := '0';
    AR_AM_O5	: out std_logic := '0';
    AR_AM_O4	: out std_logic := '0';
    AR_AM_O3	: out std_logic := '0';
    AR_AM_O2	: out std_logic := '0';
    AR_AM_O1	: out std_logic := '0';

    AR_AP_O32	: out std_logic := '0';
    AR_AP_O31	: out std_logic := '0';
    AR_AP_O30	: out std_logic := '0';
    AR_AP_O29	: out std_logic := '0';
    AR_AP_O28	: out std_logic := '0';
    AR_AP_O27	: out std_logic := '0';
    AR_AP_O26	: out std_logic := '0';
    AR_AP_O25	: out std_logic := '0';
    AR_AP_O24	: out std_logic := '0';
    AR_AP_O23	: out std_logic := '0';
    AR_AP_O22	: out std_logic := '0';
    AR_AP_O21	: out std_logic := '0';
    AR_AP_O20	: out std_logic := '0';
    AR_AP_O19	: out std_logic := '0';
    AR_AP_O18	: out std_logic := '0';
    AR_AP_O17	: out std_logic := '0';
    AR_AP_O16	: out std_logic := '0';
    AR_AP_O15	: out std_logic := '0';
    AR_AP_O14	: out std_logic := '0';
    AR_AP_O13	: out std_logic := '0';
    AR_AP_O12	: out std_logic := '0';
    AR_AP_O11	: out std_logic := '0';
    AR_AP_O10	: out std_logic := '0';
    AR_AP_O9	: out std_logic := '0';
    AR_AP_O8	: out std_logic := '0';
    AR_AP_O7	: out std_logic := '0';
    AR_AP_O6	: out std_logic := '0';
    AR_AP_O5	: out std_logic := '0';
    AR_AP_O4	: out std_logic := '0';
    AR_AP_O3	: out std_logic := '0';
    AR_AP_O2	: out std_logic := '0';
    AR_AP_O1	: out std_logic := '0';

    AR_BUM_O2	: out std_logic := '0';
    AR_BUM_O1	: out std_logic := '0';

    AR_BUP_O2	: out std_logic := '0';
    AR_BUP_O1	: out std_logic := '0';

    AR_CHM_O4	: out std_logic := '0';
    AR_CHM_O3	: out std_logic := '0';
    AR_CHM_O2	: out std_logic := '0';
    AR_CHM_O1	: out std_logic := '0';

    AR_CHP_O4	: out std_logic := '0';
    AR_CHP_O3	: out std_logic := '0';
    AR_CHP_O2	: out std_logic := '0';
    AR_CHP_O1	: out std_logic := '0';

    AR_IDM_O4	: out std_logic := '0';
    AR_IDM_O3	: out std_logic := '0';
    AR_IDM_O2	: out std_logic := '0';
    AR_IDM_O1	: out std_logic := '0';

    AR_IDP_O4	: out std_logic := '0';
    AR_IDP_O3	: out std_logic := '0';
    AR_IDP_O2	: out std_logic := '0';
    AR_IDP_O1	: out std_logic := '0';

    AR_INM_O4	: out std_logic := '0';
    AR_INM_O3	: out std_logic := '0';
    AR_INM_O2	: out std_logic := '0';
    AR_INM_O1	: out std_logic := '0';

    AR_LEM_O4	: out std_logic := '0';
    AR_LEM_O3	: out std_logic := '0';
    AR_LEM_O2	: out std_logic := '0';
    AR_LEM_O1	: out std_logic := '0';

    AR_LEP_O4	: out std_logic := '0';
    AR_LEP_O3	: out std_logic := '0';
    AR_LEP_O2	: out std_logic := '0';
    AR_LEP_O1	: out std_logic := '0';

    AR_LKM_O2	: out std_logic := '0';
    AR_LKM_O1	: out std_logic := '0';

    AR_LKP_O2	: out std_logic := '0';
    AR_LKP_O1	: out std_logic := '0';

    AR_PRM_O3	: out std_logic := '0';
    AR_PRM_O2	: out std_logic := '0';
    AR_PRM_O1	: out std_logic := '0';

    AR_PRP_O3	: out std_logic := '0';
    AR_PRP_O2	: out std_logic := '0';
    AR_PRP_O1	: out std_logic := '0';

    AR_RDY_O	: out std_logic := '0';
    AR_SHM_O	: out std_logic := '0';

    AR_SZM_O3	: out std_logic := '0';
    AR_SZM_O2	: out std_logic := '0';
    AR_SZM_O1	: out std_logic := '0';

    AR_SZP_O3	: out std_logic := '0';
    AR_SZP_O2	: out std_logic := '0';
    AR_SZP_O1	: out std_logic := '0';

    AR_VDM_O	: out std_logic := '0';
    AR_VDP_O	: out std_logic := '0';

    AW_AM_O32	: out std_logic := '0';
    AW_AM_O31	: out std_logic := '0';
    AW_AM_O30	: out std_logic := '0';
    AW_AM_O29	: out std_logic := '0';
    AW_AM_O28	: out std_logic := '0';
    AW_AM_O27	: out std_logic := '0';
    AW_AM_O26	: out std_logic := '0';
    AW_AM_O25	: out std_logic := '0';
    AW_AM_O24	: out std_logic := '0';
    AW_AM_O23	: out std_logic := '0';
    AW_AM_O22	: out std_logic := '0';
    AW_AM_O21	: out std_logic := '0';
    AW_AM_O20	: out std_logic := '0';
    AW_AM_O19	: out std_logic := '0';
    AW_AM_O18	: out std_logic := '0';
    AW_AM_O17	: out std_logic := '0';
    AW_AM_O16	: out std_logic := '0';
    AW_AM_O15	: out std_logic := '0';
    AW_AM_O14	: out std_logic := '0';
    AW_AM_O13	: out std_logic := '0';
    AW_AM_O12	: out std_logic := '0';
    AW_AM_O11	: out std_logic := '0';
    AW_AM_O10	: out std_logic := '0';
    AW_AM_O9	: out std_logic := '0';
    AW_AM_O8	: out std_logic := '0';
    AW_AM_O7	: out std_logic := '0';
    AW_AM_O6	: out std_logic := '0';
    AW_AM_O5	: out std_logic := '0';
    AW_AM_O4	: out std_logic := '0';
    AW_AM_O3	: out std_logic := '0';
    AW_AM_O2	: out std_logic := '0';
    AW_AM_O1	: out std_logic := '0';

    AW_AP_O32	: out std_logic := '0';
    AW_AP_O31	: out std_logic := '0';
    AW_AP_O30	: out std_logic := '0';
    AW_AP_O29	: out std_logic := '0';
    AW_AP_O28	: out std_logic := '0';
    AW_AP_O27	: out std_logic := '0';
    AW_AP_O26	: out std_logic := '0';
    AW_AP_O25	: out std_logic := '0';
    AW_AP_O24	: out std_logic := '0';
    AW_AP_O23	: out std_logic := '0';
    AW_AP_O22	: out std_logic := '0';
    AW_AP_O21	: out std_logic := '0';
    AW_AP_O20	: out std_logic := '0';
    AW_AP_O19	: out std_logic := '0';
    AW_AP_O18	: out std_logic := '0';
    AW_AP_O17	: out std_logic := '0';
    AW_AP_O16	: out std_logic := '0';
    AW_AP_O15	: out std_logic := '0';
    AW_AP_O14	: out std_logic := '0';
    AW_AP_O13	: out std_logic := '0';
    AW_AP_O12	: out std_logic := '0';
    AW_AP_O11	: out std_logic := '0';
    AW_AP_O10	: out std_logic := '0';
    AW_AP_O9	: out std_logic := '0';
    AW_AP_O8	: out std_logic := '0';
    AW_AP_O7	: out std_logic := '0';
    AW_AP_O6	: out std_logic := '0';
    AW_AP_O5	: out std_logic := '0';
    AW_AP_O4	: out std_logic := '0';
    AW_AP_O3	: out std_logic := '0';
    AW_AP_O2	: out std_logic := '0';
    AW_AP_O1	: out std_logic := '0';

    AW_BUM_O2	: out std_logic := '0';
    AW_BUM_O1	: out std_logic := '0';

    AW_BUP_O2	: out std_logic := '0';
    AW_BUP_O1	: out std_logic := '0';

    AW_CHM_O4	: out std_logic := '0';
    AW_CHM_O3	: out std_logic := '0';
    AW_CHM_O2	: out std_logic := '0';
    AW_CHM_O1	: out std_logic := '0';

    AW_CHP_O4	: out std_logic := '0';
    AW_CHP_O3	: out std_logic := '0';
    AW_CHP_O2	: out std_logic := '0';
    AW_CHP_O1	: out std_logic := '0';

    AW_IDM_O4	: out std_logic := '0';
    AW_IDM_O3	: out std_logic := '0';
    AW_IDM_O2	: out std_logic := '0';
    AW_IDM_O1	: out std_logic := '0';

    AW_IDP_O4	: out std_logic := '0';
    AW_IDP_O3	: out std_logic := '0';
    AW_IDP_O2	: out std_logic := '0';
    AW_IDP_O1	: out std_logic := '0';

    AW_INM_O4	: out std_logic := '0';
    AW_INM_O3	: out std_logic := '0';
    AW_INM_O2	: out std_logic := '0';
    AW_INM_O1	: out std_logic := '0';

    AW_LEM_O4	: out std_logic := '0';
    AW_LEM_O3	: out std_logic := '0';
    AW_LEM_O2	: out std_logic := '0';
    AW_LEM_O1	: out std_logic := '0';

    AW_LEP_O4	: out std_logic := '0';
    AW_LEP_O3	: out std_logic := '0';
    AW_LEP_O2	: out std_logic := '0';
    AW_LEP_O1	: out std_logic := '0';

    AW_LKM_O2	: out std_logic := '0';
    AW_LKM_O1	: out std_logic := '0';

    AW_LKP_O2	: out std_logic := '0';
    AW_LKP_O1	: out std_logic := '0';

    AW_PRM_O3	: out std_logic := '0';
    AW_PRM_O2	: out std_logic := '0';
    AW_PRM_O1	: out std_logic := '0';

    AW_PRP_O3	: out std_logic := '0';
    AW_PRP_O2	: out std_logic := '0';
    AW_PRP_O1	: out std_logic := '0';

    AW_RDY_O	: out std_logic := '0';
    AW_SHM_O	: out std_logic := '0';

    AW_SZM_O3	: out std_logic := '0';
    AW_SZM_O2	: out std_logic := '0';
    AW_SZM_O1	: out std_logic := '0';

    AW_SZP_O3	: out std_logic := '0';
    AW_SZP_O2	: out std_logic := '0';
    AW_SZP_O1	: out std_logic := '0';

    AW_VDM_O	: out std_logic := '0';
    AW_VDP_O	: out std_logic := '0';

    B_IDS_O8	: out std_logic := '0';
    B_IDS_O7	: out std_logic := '0';
    B_IDS_O6	: out std_logic := '0';
    B_IDS_O5	: out std_logic := '0';
    B_IDS_O4	: out std_logic := '0';
    B_IDS_O3	: out std_logic := '0';
    B_IDS_O2	: out std_logic := '0';
    B_IDS_O1	: out std_logic := '0';

    B_RDYM_O	: out std_logic := '0';
    B_RDYP_O	: out std_logic := '0';

    B_RSP_O2	: out std_logic := '0';
    B_RSP_O1	: out std_logic := '0';

    B_VD_O	: out std_logic := '0';

--    CAL_O5        : out std_logic; --  calibration         5   [0:4]
--    CAL_O4        : out std_logic; --  calibration         5   [0:4]
--    CAL_O3        : out std_logic; --  calibration         5   [0:4]
--    CAL_O2        : out std_logic; --  calibration         5   [0:4]
--    CAL_O1        : out std_logic; --  calibration         5   [0:4]

    CDB_PW_O	: out std_logic := '0';
    CDB_RS_O	: out std_logic := '0';
--    CK_DR_O       : out std_logic; --  clock_dr            1
    COM_RX_O	: out std_logic := '0';
    COM_TX_O	: out std_logic := '0';
    CS_PW_O	: out std_logic := '0';
    DB_ACK_O	: out std_logic := '0';
    DB_NPD_O	: out std_logic := '0';
    DB_RS_O	: out std_logic := '0';

    DFTS_O8	: out std_logic := '0';
    DFTS_O7	: out std_logic := '0';
    DFTS_O6	: out std_logic := '0';
    DFTS_O5	: out std_logic := '0';
    DFTS_O4	: out std_logic := '0';
    DFTS_O3	: out std_logic := '0';
    DFTS_O2	: out std_logic := '0';
    DFTS_O1	: out std_logic := '0';

    ET_ASC_O8	: out std_logic := '0';
    ET_ASC_O7	: out std_logic := '0';
    ET_ASC_O6	: out std_logic := '0';
    ET_ASC_O5	: out std_logic := '0';
    ET_ASC_O4	: out std_logic := '0';
    ET_ASC_O3	: out std_logic := '0';
    ET_ASC_O2	: out std_logic := '0';
    ET_ASC_O1	: out std_logic := '0';

    ET_E_O	: out std_logic := '0';

    ET_EXT_O2	: out std_logic := '0';
    ET_EXT_O1	: out std_logic := '0';

    EVENT_O	: out std_logic := '0';
    FP_DZC_O	: out std_logic := '0';
    FP_IDC_O	: out std_logic := '0';
    FP_IOC_O	: out std_logic := '0';
    FP_IXC_O	: out std_logic := '0';
    FP_OFC_O	: out std_logic := '0';
    FP_UFC_O	: out std_logic := '0';
    JTAG_O	: out std_logic := '0';
--    LBK_E_O       : out std_logic; --  loopback_en         1
--    LBK_MX_O      : out std_logic; --  loopback_mux        1

--    MODE1_O2      : out std_logic; --  mode1               3   [0:2]
--    MODE1_O1      : out std_logic; --  mode1               3   [0:2]

--    MODE2_O2      : out std_logic; --  mode2               3   [0:2]
--    MODE2_O1      : out std_logic; --  mode2               3   [0:2]

--    MODE3_O2      : out std_logic; --  mode3               3   [0:2]
--    MODE3_O1      : out std_logic; --  mode3               3   [0:2]

    N_CKST_O	: out std_logic := '0';
    N_PMU_O	: out std_logic := '0';
    N_TDO_O	: out std_logic := '0';
    N_VFIQ_O	: out std_logic := '0';
    N_VIRQ_O	: out std_logic := '0';
    N_VRST_O	: out std_logic := '0';
    N_EPST_O	: out std_logic := '0';
    N_IPST_O	: out std_logic := '0';

    P_RD_O32	: out std_logic := '0';
    P_RD_O31	: out std_logic := '0';
    P_RD_O30	: out std_logic := '0';
    P_RD_O29	: out std_logic := '0';
    P_RD_O28	: out std_logic := '0';
    P_RD_O27	: out std_logic := '0';
    P_RD_O26	: out std_logic := '0';
    P_RD_O25	: out std_logic := '0';
    P_RD_O24	: out std_logic := '0';
    P_RD_O23	: out std_logic := '0';
    P_RD_O22	: out std_logic := '0';
    P_RD_O21	: out std_logic := '0';
    P_RD_O20	: out std_logic := '0';
    P_RD_O19	: out std_logic := '0';
    P_RD_O18	: out std_logic := '0';
    P_RD_O17	: out std_logic := '0';
    P_RD_O16	: out std_logic := '0';
    P_RD_O15	: out std_logic := '0';
    P_RD_O14	: out std_logic := '0';
    P_RD_O13	: out std_logic := '0';
    P_RD_O12	: out std_logic := '0';
    P_RD_O11	: out std_logic := '0';
    P_RD_O10	: out std_logic := '0';
    P_RD_O9	: out std_logic := '0';
    P_RD_O8	: out std_logic := '0';
    P_RD_O7	: out std_logic := '0';
    P_RD_O6	: out std_logic := '0';
    P_RD_O5	: out std_logic := '0';
    P_RD_O4	: out std_logic := '0';
    P_RD_O3	: out std_logic := '0';
    P_RD_O2	: out std_logic := '0';
    P_RD_O1	: out std_logic := '0';

    P_RDY_O	: out std_logic := '0';
    P_VER_O	: out std_logic := '0';

    RD_O64	: out std_logic := '0';
    RD_O63	: out std_logic := '0';
    RD_O62	: out std_logic := '0';
    RD_O61	: out std_logic := '0';
    RD_O60	: out std_logic := '0';
    RD_O59	: out std_logic := '0';
    RD_O58	: out std_logic := '0';
    RD_O57	: out std_logic := '0';
    RD_O56	: out std_logic := '0';
    RD_O55	: out std_logic := '0';
    RD_O54	: out std_logic := '0';
    RD_O53	: out std_logic := '0';
    RD_O52	: out std_logic := '0';
    RD_O51	: out std_logic := '0';
    RD_O50	: out std_logic := '0';
    RD_O49	: out std_logic := '0';
    RD_O48	: out std_logic := '0';
    RD_O47	: out std_logic := '0';
    RD_O46	: out std_logic := '0';
    RD_O45	: out std_logic := '0';
    RD_O44	: out std_logic := '0';
    RD_O43	: out std_logic := '0';
    RD_O42	: out std_logic := '0';
    RD_O41	: out std_logic := '0';
    RD_O40	: out std_logic := '0';
    RD_O39	: out std_logic := '0';
    RD_O38	: out std_logic := '0';
    RD_O37	: out std_logic := '0';
    RD_O36	: out std_logic := '0';
    RD_O35	: out std_logic := '0';
    RD_O34	: out std_logic := '0';
    RD_O33	: out std_logic := '0';
    RD_O32	: out std_logic := '0';
    RD_O31	: out std_logic := '0';
    RD_O30	: out std_logic := '0';
    RD_O29	: out std_logic := '0';
    RD_O28	: out std_logic := '0';
    RD_O27	: out std_logic := '0';
    RD_O26	: out std_logic := '0';
    RD_O25	: out std_logic := '0';
    RD_O24	: out std_logic := '0';
    RD_O23	: out std_logic := '0';
    RD_O22	: out std_logic := '0';
    RD_O21	: out std_logic := '0';
    RD_O20	: out std_logic := '0';
    RD_O19	: out std_logic := '0';
    RD_O18	: out std_logic := '0';
    RD_O17	: out std_logic := '0';
    RD_O16	: out std_logic := '0';
    RD_O15	: out std_logic := '0';
    RD_O14	: out std_logic := '0';
    RD_O13	: out std_logic := '0';
    RD_O12	: out std_logic := '0';
    RD_O11	: out std_logic := '0';
    RD_O10	: out std_logic := '0';
    RD_O9	: out std_logic := '0';
    RD_O8	: out std_logic := '0';
    RD_O7	: out std_logic := '0';
    RD_O6	: out std_logic := '0';
    RD_O5	: out std_logic := '0';
    RD_O4	: out std_logic := '0';
    RD_O3	: out std_logic := '0';
    RD_O2	: out std_logic := '0';
    RD_O1	: out std_logic := '0';

--    RDY_O3        : out std_logic; --  ready               3   [0:2]
--    RDY_O2        : out std_logic; --  ready               3   [0:2]
--    RDY_O1        : out std_logic; --  ready               3   [0:2]

    R_IDS_O8	: out std_logic := '0';
    R_IDS_O7	: out std_logic := '0';
    R_IDS_O6	: out std_logic := '0';
    R_IDS_O5	: out std_logic := '0';
    R_IDS_O4	: out std_logic := '0';
    R_IDS_O3	: out std_logic := '0';
    R_IDS_O2	: out std_logic := '0';
    R_IDS_O1	: out std_logic := '0';

    R_LST_O	: out std_logic := '0';
    R_RDYM_O	: out std_logic := '0';
    R_RDYP_O	: out std_logic := '0';

    R_RSP_O2	: out std_logic := '0';
    R_RSP_O1	: out std_logic := '0';

    R_VD_O	: out std_logic := '0';
--    SCAN_E_O      : out std_logic; --  scan_en             1
--    SHF_DR_O      : out std_logic; --  shift_dr            1
--    SHOUT_O       : out std_logic; --  shout               1
    SWDO_O	: out std_logic := '0';
    SWDO_E_O	: out std_logic := '0';
    TDO_O	: out std_logic := '0';
--    TEST_E_O      : out std_logic; --  test_en             1
    T_CK_O	: out std_logic := '0';
    T_CTL_O	: out std_logic := '0';

    T_DATA_O32	: out std_logic := '0';
    T_DATA_O31	: out std_logic := '0';
    T_DATA_O30	: out std_logic := '0';
    T_DATA_O29	: out std_logic := '0';
    T_DATA_O28	: out std_logic := '0';
    T_DATA_O27	: out std_logic := '0';
    T_DATA_O26	: out std_logic := '0';
    T_DATA_O25	: out std_logic := '0';
    T_DATA_O24	: out std_logic := '0';
    T_DATA_O23	: out std_logic := '0';
    T_DATA_O22	: out std_logic := '0';
    T_DATA_O21	: out std_logic := '0';
    T_DATA_O20	: out std_logic := '0';
    T_DATA_O19	: out std_logic := '0';
    T_DATA_O18	: out std_logic := '0';
    T_DATA_O17	: out std_logic := '0';
    T_DATA_O16	: out std_logic := '0';
    T_DATA_O15	: out std_logic := '0';
    T_DATA_O14	: out std_logic := '0';
    T_DATA_O13	: out std_logic := '0';
    T_DATA_O12	: out std_logic := '0';
    T_DATA_O11	: out std_logic := '0';
    T_DATA_O10	: out std_logic := '0';
    T_DATA_O9	: out std_logic := '0';
    T_DATA_O8	: out std_logic := '0';
    T_DATA_O7	: out std_logic := '0';
    T_DATA_O6	: out std_logic := '0';
    T_DATA_O5	: out std_logic := '0';
    T_DATA_O4	: out std_logic := '0';
    T_DATA_O3	: out std_logic := '0';
    T_DATA_O2	: out std_logic := '0';
    T_DATA_O1	: out std_logic := '0';

--    UPD_DR_O      : out std_logic; --  update_dr           1

    W_DM_O64	: out std_logic := '0';
    W_DM_O63	: out std_logic := '0';
    W_DM_O62	: out std_logic := '0';
    W_DM_O61	: out std_logic := '0';
    W_DM_O60	: out std_logic := '0';
    W_DM_O59	: out std_logic := '0';
    W_DM_O58	: out std_logic := '0';
    W_DM_O57	: out std_logic := '0';
    W_DM_O56	: out std_logic := '0';
    W_DM_O55	: out std_logic := '0';
    W_DM_O54	: out std_logic := '0';
    W_DM_O53	: out std_logic := '0';
    W_DM_O52	: out std_logic := '0';
    W_DM_O51	: out std_logic := '0';
    W_DM_O50	: out std_logic := '0';
    W_DM_O49	: out std_logic := '0';
    W_DM_O48	: out std_logic := '0';
    W_DM_O47	: out std_logic := '0';
    W_DM_O46	: out std_logic := '0';
    W_DM_O45	: out std_logic := '0';
    W_DM_O44	: out std_logic := '0';
    W_DM_O43	: out std_logic := '0';
    W_DM_O42	: out std_logic := '0';
    W_DM_O41	: out std_logic := '0';
    W_DM_O40	: out std_logic := '0';
    W_DM_O39	: out std_logic := '0';
    W_DM_O38	: out std_logic := '0';
    W_DM_O37	: out std_logic := '0';
    W_DM_O36	: out std_logic := '0';
    W_DM_O35	: out std_logic := '0';
    W_DM_O34	: out std_logic := '0';
    W_DM_O33	: out std_logic := '0';
    W_DM_O32	: out std_logic := '0';
    W_DM_O31	: out std_logic := '0';
    W_DM_O30	: out std_logic := '0';
    W_DM_O29	: out std_logic := '0';
    W_DM_O28	: out std_logic := '0';
    W_DM_O27	: out std_logic := '0';
    W_DM_O26	: out std_logic := '0';
    W_DM_O25	: out std_logic := '0';
    W_DM_O24	: out std_logic := '0';
    W_DM_O23	: out std_logic := '0';
    W_DM_O22	: out std_logic := '0';
    W_DM_O21	: out std_logic := '0';
    W_DM_O20	: out std_logic := '0';
    W_DM_O19	: out std_logic := '0';
    W_DM_O18	: out std_logic := '0';
    W_DM_O17	: out std_logic := '0';
    W_DM_O16	: out std_logic := '0';
    W_DM_O15	: out std_logic := '0';
    W_DM_O14	: out std_logic := '0';
    W_DM_O13	: out std_logic := '0';
    W_DM_O12	: out std_logic := '0';
    W_DM_O11	: out std_logic := '0';
    W_DM_O10	: out std_logic := '0';
    W_DM_O9	: out std_logic := '0';
    W_DM_O8	: out std_logic := '0';
    W_DM_O7	: out std_logic := '0';
    W_DM_O6	: out std_logic := '0';
    W_DM_O5	: out std_logic := '0';
    W_DM_O4	: out std_logic := '0';
    W_DM_O3	: out std_logic := '0';
    W_DM_O2	: out std_logic := '0';
    W_DM_O1	: out std_logic := '0';

    W_DP_O32	: out std_logic := '0';
    W_DP_O31	: out std_logic := '0';
    W_DP_O30	: out std_logic := '0';
    W_DP_O29	: out std_logic := '0';
    W_DP_O28	: out std_logic := '0';
    W_DP_O27	: out std_logic := '0';
    W_DP_O26	: out std_logic := '0';
    W_DP_O25	: out std_logic := '0';
    W_DP_O24	: out std_logic := '0';
    W_DP_O23	: out std_logic := '0';
    W_DP_O22	: out std_logic := '0';
    W_DP_O21	: out std_logic := '0';
    W_DP_O20	: out std_logic := '0';
    W_DP_O19	: out std_logic := '0';
    W_DP_O18	: out std_logic := '0';
    W_DP_O17	: out std_logic := '0';
    W_DP_O16	: out std_logic := '0';
    W_DP_O15	: out std_logic := '0';
    W_DP_O14	: out std_logic := '0';
    W_DP_O13	: out std_logic := '0';
    W_DP_O12	: out std_logic := '0';
    W_DP_O11	: out std_logic := '0';
    W_DP_O10	: out std_logic := '0';
    W_DP_O9	: out std_logic := '0';
    W_DP_O8	: out std_logic := '0';
    W_DP_O7	: out std_logic := '0';
    W_DP_O6	: out std_logic := '0';
    W_DP_O5	: out std_logic := '0';
    W_DP_O4	: out std_logic := '0';
    W_DP_O3	: out std_logic := '0';
    W_DP_O2	: out std_logic := '0';
    W_DP_O1	: out std_logic := '0';

    W_IDM_O4	: out std_logic := '0';
    W_IDM_O3	: out std_logic := '0';
    W_IDM_O2	: out std_logic := '0';
    W_IDM_O1	: out std_logic := '0';

    W_IDP_O4	: out std_logic := '0';
    W_IDP_O3	: out std_logic := '0';
    W_IDP_O2	: out std_logic := '0';
    W_IDP_O1	: out std_logic := '0';

    W_LSTM_O	: out std_logic := '0';
    W_LSTP_O	: out std_logic := '0';
    W_RDY_O	: out std_logic := '0';

    W_SBM_O8	: out std_logic := '0';
    W_SBM_O7	: out std_logic := '0';
    W_SBM_O6	: out std_logic := '0';
    W_SBM_O5	: out std_logic := '0';
    W_SBM_O4	: out std_logic := '0';
    W_SBM_O3	: out std_logic := '0';
    W_SBM_O2	: out std_logic := '0';
    W_SBM_O1	: out std_logic := '0';

    W_SBP_O4	: out std_logic := '0';
    W_SBP_O3	: out std_logic := '0';
    W_SBP_O2	: out std_logic := '0';
    W_SBP_O1	: out std_logic := '0';

    W_VDM_O	: out std_logic := '0';
    W_VDP_O	: out std_logic := '0'
);
end component NX_R5_L;

component NX_R5_L_WRAP is
port (
            ------------------------------------------------------------------------
            -- CORTEXR5 PRIMARY INPUTS AND OUTPUTS
            ------------------------------------------------------------------------  
            ------------------------------------------------------------------------
            -- Global
            ------------------------------------------------------------------------
    CLKIN	: in std_logic := '0';
    nRESET0	: in std_logic := '0';
    nSYSPORESET	: in std_logic := '0';
    nCPUHALT0	: in std_logic := '0';
    DBGNOCLKSTOP	: in std_logic := '0';
    nCLKSTOPPED0	: out std_logic := '0';
    nWFEPIPESTOPPED0	: out std_logic := '0';
    nWFIPIPESTOPPED0	: out std_logic := '0';
    EVENTI0	: in std_logic := '0';
    EVENTO0	: out std_logic := '0';
            ------------------------------------------------------------------------
            -- Configuration signals
            ------------------------------------------------------------------------
    VINITHI0	: in std_logic := '0';
    CFGEE	: in std_logic := '0';
    CFGIE	: in std_logic := '0';
    INITRAMA0	: in std_logic := '0';
    LOCZRAMA0	: in std_logic := '0';
    TEINIT	: in std_logic := '0';
    CFGNMFI0	: in std_logic := '0';
    PARECCENRAM0	: in std_logic := '0';
    PARITYLEVEL	: in std_logic := '0';
    ERRENRAM0	: in std_logic := '0';
    GROUPID	: in std_logic_vector(3 downto 0) := (others => '0');
    INITPPX0	: in std_logic := '0';
    PPXBASE0	: in std_logic_vector(19 downto 0) := (others => '0');
    PPXSIZE0	: in std_logic_vector(4 downto 0) := (others => '0');
    PPVBASE0	: in std_logic_vector(19 downto 0) := (others => '0');
    PPVSIZE0	: in std_logic_vector(4 downto 0) := (others => '0');
            ------------------------------------------------------------------------
            -- Interrupt signals
            ------------------------------------------------------------------------
    nFIQ0	: in std_logic := '0';
    nIRQ0	: in std_logic := '0';
    nPMUIRQ0	: out std_logic := '0';
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Master Port
            ------------------------------------------------------------------------
    ACLKENM0	: in std_logic := '0';
            -- Write Address Channel
    AWADDRM0	: out std_logic_vector(31 downto 0) := (others => '0');
    AWBURSTM0	: out std_logic_vector(1 downto 0) := (others => '0');
    AWCACHEM0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWIDM0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWLENM0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWLOCKM0	: out std_logic_vector(1 downto 0) := (others => '0');
    AWPROTM0	: out std_logic_vector(2 downto 0) := (others => '0');
    AWREADYM0	: in std_logic := '0';
    AWSIZEM0	: out std_logic_vector(2 downto 0) := (others => '0');
    AWINNERM0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWSHAREM0	: out std_logic := '0';
    AWVALIDM0	: out std_logic := '0';
            -- Write Data Channel
    WDATAM0	: out std_logic_vector(63 downto 0) := (others => '0');
    WIDM0	: out std_logic_vector(3 downto 0) := (others => '0');
    WLASTM0	: out std_logic := '0';
    WREADYM0	: in std_logic := '0';
    WSTRBM0	: out std_logic_vector(7 downto 0) := (others => '0');
    WVALIDM0	: out std_logic := '0';
            -- Write response channel
    BIDM0	: in std_logic_vector(3 downto 0) := (others => '0');
    BREADYM0	: out std_logic := '0';
    BRESPM0	: in std_logic_vector(1 downto 0) := (others => '0');
    BVALIDM0	: in std_logic := '0';
            -- Read Address Channel
    ARADDRM0	: out std_logic_vector(31 downto 0) := (others => '0');
    ARBURSTM0	: out std_logic_vector(1 downto 0) := (others => '0');
    ARCACHEM0	: out std_logic_vector(3 downto 0) := (others => '0');
    ARIDM0	: out std_logic_vector(3 downto 0) := (others => '0');
    ARLENM0	: out std_logic_vector(3 downto 0) := (others => '0');
    ARLOCKM0	: out std_logic_vector(1 downto 0) := (others => '0');
    ARPROTM0	: out std_logic_vector(2 downto 0) := (others => '0');
    ARREADYM0	: in std_logic := '0';
    ARSIZEM0	: out std_logic_vector(2 downto 0) := (others => '0');
    ARINNERM0	: out std_logic_vector(3 downto 0) := (others => '0');
    ARSHAREM0	: out std_logic := '0';
    ARVALIDM0	: out std_logic := '0';
            -- Read Data Channel
    RDATAM0	: in std_logic_vector(63 downto 0) := (others => '0');
    RIDM0	: in std_logic_vector(3 downto 0) := (others => '0');
    RLASTM0	: in std_logic := '0';
    RREADYM0	: out std_logic := '0';
    RRESPM0	: in std_logic_vector(1 downto 0) := (others => '0');
    RVALIDM0	: in std_logic := '0';
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Slave Port
            ------------------------------------------------------------------------
    ACLKENS0	: in std_logic := '0';
            -- Write Address Channel
    AWADDRS0	: in std_logic_vector(31 downto 0) := (others => '0');
    AWBURSTS0	: in std_logic_vector(1 downto 0) := (others => '0');
    AWCACHES0	: in std_logic_vector(3 downto 0) := (others => '0');

    AWIDS0	: in std_logic_vector(7 downto 0) := (others => '0');
    AWLENS0	: in std_logic_vector(3 downto 0) := (others => '0');
    AWLOCKS0	: in std_logic_vector(1 downto 0) := (others => '0');
    AWPROTS0	: in std_logic_vector(2 downto 0) := (others => '0');
    AWREADYS0	: out std_logic := '0';
    AWSIZES0	: in std_logic_vector(2 downto 0) := (others => '0');
    AWVALIDS0	: in std_logic := '0';
            -- Write Data Channel
    WDATAS0	: in std_logic_vector(63 downto 0) := (others => '0');
    WIDS0	: in std_logic_vector(7 downto 0) := (others => '0');
    WLASTS0	: in std_logic := '0';
    WREADYS0	: out std_logic := '0';
    WSTRBS0	: in std_logic_vector(7 downto 0) := (others => '0');
    WVALIDS0	: in std_logic := '0';
            -- Write response channel
    BIDS0	: out std_logic_vector(7 downto 0) := (others => '0');
    BREADYS0	: in std_logic := '0';
    BRESPS0	: out std_logic_vector(1 downto 0) := (others => '0');
    BVALIDS0	: out std_logic := '0';
            -- Read Address Channel
    ARADDRS0	: in std_logic_vector(31 downto 0) := (others => '0');
    ARBURSTS0	: in std_logic_vector(1 downto 0) := (others => '0');
    ARCACHES0	: in std_logic_vector(3 downto 0) := (others => '0');
    ARIDS0	: in std_logic_vector(7 downto 0) := (others => '0');
    ARLENS0	: in std_logic_vector(3 downto 0) := (others => '0');
    ARLOCKS0	: in std_logic_vector(1 downto 0) := (others => '0');
    ARPROTS0	: in std_logic_vector(2 downto 0) := (others => '0');
    ARREADYS0	: out std_logic := '0';
    ARSIZES0	: in std_logic_vector(2 downto 0) := (others => '0');

    ARVALIDS0	: in std_logic := '0';
            -- Read Data Channel
    RDATAS0	: out std_logic_vector(63 downto 0) := (others => '0');
    RIDS0	: out std_logic_vector(7 downto 0) := (others => '0');
    RLASTS0	: out std_logic := '0';
    RREADYS0	: in std_logic := '0';
    RRESPS0	: out std_logic_vector(1 downto 0) := (others => '0');
    RVALIDS0	: out std_logic := '0';
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Peripheral Port
            ------------------------------------------------------------------------
    ACLKENP0	: in std_logic := '0';
            -- Write Address Channel
    AWIDP0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWADDRP0	: out std_logic_vector(31 downto 0) := (others => '0');
    AWLENP0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWSIZEP0	: out std_logic_vector(2 downto 0) := (others => '0');
    AWBURSTP0	: out std_logic_vector(1 downto 0) := (others => '0');
    AWLOCKP0	: out std_logic_vector(1 downto 0) := (others => '0');
    AWCACHEP0	: out std_logic_vector(3 downto 0) := (others => '0');
    AWPROTP0	: out std_logic_vector(2 downto 0) := (others => '0');
    AWVALIDP0	: out std_logic := '0';
    AWREADYP0	: in std_logic := '0';
            -- Write Data Channel
    WIDP0	: out std_logic_vector(3 downto 0) := (others => '0');
    WDATAP0	: out std_logic_vector(31 downto 0) := (others => '0');
    WSTRBP0	: out std_logic_vector(3 downto 0) := (others => '0');
    WLASTP0	: out std_logic := '0';
    WVALIDP0	: out std_logic := '0';
    WREADYP0	: in std_logic := '0';
            -- Write response channel
    BIDP0	: in std_logic_vector(3 downto 0) := (others => '0');
    BRESPP0	: in std_logic_vector(1 downto 0) := (others => '0');
    BVALIDP0	: in std_logic := '0';
    BREADYP0	: out std_logic := '0';
            -- Read Address Channel
            ARIDP0       : out std_logic_vector (3 downto 0);          
            ARADDRP0     : out std_logic_vector (31 downto 0);          
            ARLENP0      : out std_logic_vector (3 downto 0);          
            ARSIZEP0     : out std_logic_vector (2 downto 0);          
            ARBURSTP0    : out std_logic_vector (1 downto 0);          
            ARLOCKP0     : out std_logic_vector (1 downto 0);          
            ARCACHEP0    : out std_logic_vector (3 downto 0);          
            ARPROTP0     : out std_logic_vector (2 downto 0);          
    ARVALIDP0	: out std_logic := '0';
    ARREADYP0	: in std_logic := '0';
            -- Reainata Channel
    RIDP0	: in std_logic_vector(3 downto 0) := (others => '0');
    RDATAP0	: in std_logic_vector(31 downto 0) := (others => '0');
    RRESPP0	: in std_logic_vector(1 downto 0) := (others => '0');
    RLASTP0	: in std_logic := '0';
    RVALIDP0	: in std_logic := '0';
    RREADYP0	: out std_logic := '0';
       
            -- Debug Miscellaneous
    DBGEN0	: in std_logic := '0';
    NIDEN0	: in std_logic := '0';
    EDBGRQ0	: in std_logic := '0';
    DBGACK0	: out std_logic := '0';
    DBGRSTREQ0	: out std_logic := '0';

    COMMRX0	: out std_logic := '0';
    COMMTX0	: out std_logic := '0';

    DBGNOPWRDWN	: out std_logic := '0';
    DBGROMADDR	: in std_logic_vector(19 downto 0) := (others => '0');
    DBGROMADDRV	: in std_logic := '0';
    DBGSELFADDR0	: in std_logic_vector(19 downto 0) := (others => '0');
    DBGSELFADDRV0	: in std_logic := '0';
            ------------------------------------------------------------------------
            -- ETM Interface
            ------------------------------------------------------------------------
    nETMPORESET	: in std_logic := '0';
    ETMASICCTL0	: out std_logic_vector(7 downto 0) := (others => '0');
    ETMEN0	: out std_logic := '0';
    ETMEXTOUT0	: out std_logic_vector(1 downto 0) := (others => '0');
            ------------------------------------------------------------------------
            -- Validation
            ------------------------------------------------------------------------
    nVALIRQ0	: out std_logic := '0';
    nVALFIQ0	: out std_logic := '0';
    nVALRESET0	: out std_logic := '0';
       
            ------------------------------------------------------------------------
            -- FPU
            ------------------------------------------------------------------------
    FPIXC0	: out std_logic := '0';
    FPOFC0	: out std_logic := '0';
    FPUFC0	: out std_logic := '0';
    FPIOC0	: out std_logic := '0';
    FPDZC0	: out std_logic := '0';
    FPIDC0	: out std_logic := '0';
            ------------------------------------------------------------------------
            -- Coresight TPIU-Lite
            ------------------------------------------------------------------------
            ------------------------------------------------------------------------
            -- ATB Port
            ------------------------------------------------------------------------
    ATRESETn	: in std_logic := '0';
            ------------------------------------------------------------------------
            -- Trace Out Port
            ------------------------------------------------------------------------
    TRACECLK	: out std_logic := '0';
    TRACEDATA	: out std_logic_vector(31 downto 0) := (others => '0');
    TRACECTL	: out std_logic := '0';
            ------------------------------------------------------------------------
            -- Coresight DAP-Lite
            ------------------------------------------------------------------------
            ------------------------------------------------------------------------
            -- CoreSight DAP Ports
            ------------------------------------------------------------------------    
    PCLKSYS	: in std_logic := '0';
    PCLKENSYS	: in std_logic := '0';
    PRESETSYSn	: in std_logic := '0';
    PADDRSYS	: in std_logic_vector(28 downto 0) := (others => '0');
    PENABLESYS	: in std_logic := '0';
    PRDATASYS	: out std_logic_vector(31 downto 0) := (others => '0');
    PREADYSYS	: out std_logic := '0';
    PSELSYS	: in std_logic := '0';
    PSLVERRSYS	: out std_logic := '0';
    PWDATASYS	: in std_logic_vector(31 downto 0) := (others => '0');
    PWRITESYS	: in std_logic := '0';
       
    CDBGPWRUPACK	: in std_logic := '0';
    CDBGPWRUPREQ	: out std_logic := '0';
    CDBGRSTACK	: in std_logic := '0';
    CDBGRSTREQ	: out std_logic := '0';
    CSYSPWRUPACK	: in std_logic := '0';
    CSYSPWRUPREQ	: out std_logic := '0';
    DEVICEEN	: in std_logic := '0';
    JTAGNSW	: out std_logic := '0';
    nPOTRST	: in std_logic := '0';
    nTDOEN	: out std_logic := '0';
    nTRST	: in std_logic := '0';
    SWCLKTCK	: in std_logic := '0';
    SWDITMS	: in std_logic := '0';
    SWDO	: out std_logic := '0';
    SWDOEN	: out std_logic := '0';
    TDI	: in std_logic := '0';
    TDO	: out std_logic := '0'

);
end component NX_R5_L_WRAP;

component NX_RB is
generic (
    -- input : EI to FO
    inputClk      : bit_vector( 1 downto 0) := B"00"; -- 00 = CK1, 01 = CK2, 10 = CK3 and 11 = CK4
    inputBypass   : bit_vector(23 downto 0) := B"000000000000000000000000"; -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    inputContext  : string := ""; -- input context initialization
    -- output : FI to EO
    outputClk     : bit_vector( 1 downto 0) := B"00"; -- 00 = CK1, 01 = CK2, 10 = CK3 and 11 = CK4
    outputBypass  : bit_vector(23 downto 0) := B"000000000000000000000000";  -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    outputContext : string := "" -- output context initialization
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    CK3	: in std_logic := '0';
    CK4	: in std_logic := '0';
    EI1	: in std_logic := '0';
    EI2	: in std_logic := '0';
    EI3	: in std_logic := '0';
    EI4	: in std_logic := '0';
    EI5	: in std_logic := '0';
    EI6	: in std_logic := '0';
    EI7	: in std_logic := '0';
    EI8	: in std_logic := '0';
    EI9	: in std_logic := '0';
    EI10	: in std_logic := '0';
    EI11	: in std_logic := '0';
    EI12	: in std_logic := '0';
    EI13	: in std_logic := '0';
    EI14	: in std_logic := '0';
    EI15	: in std_logic := '0';
    EI16	: in std_logic := '0';
    EI17	: in std_logic := '0';
    EI18	: in std_logic := '0';
    EI19	: in std_logic := '0';
    EI20	: in std_logic := '0';
    EI21	: in std_logic := '0';
    EI22	: in std_logic := '0';
    EI23	: in std_logic := '0';
    EI24	: in std_logic := '0';
    EI25	: in std_logic := '0';
    EI26	: in std_logic := '0';
    EI27	: in std_logic := '0';
    EI28	: in std_logic := '0';
    EI29	: in std_logic := '0';
    EI30	: in std_logic := '0';
    EI31	: in std_logic := '0';
    EI32	: in std_logic := '0';
    EI33	: in std_logic := '0';
    EI34	: in std_logic := '0';
    EI35	: in std_logic := '0';
    EI36	: in std_logic := '0';
    EI37	: in std_logic := '0';
    EI38	: in std_logic := '0';
    EI39	: in std_logic := '0';
    EI40	: in std_logic := '0';
    EI41	: in std_logic := '0';
    EI42	: in std_logic := '0';
    EI43	: in std_logic := '0';
    EI44	: in std_logic := '0';
    EI45	: in std_logic := '0';
    EI46	: in std_logic := '0';
    EI47	: in std_logic := '0';
    EI48	: in std_logic := '0';
    EI49	: in std_logic := '0';
    EI50	: in std_logic := '0';
    EI51	: in std_logic := '0';
    EI52	: in std_logic := '0';
    EI53	: in std_logic := '0';
    EI54	: in std_logic := '0';
    EI55	: in std_logic := '0';
    EI56	: in std_logic := '0';
    EI57	: in std_logic := '0';
    EI58	: in std_logic := '0';
    EI59	: in std_logic := '0';
    EI60	: in std_logic := '0';
    EI61	: in std_logic := '0';
    EI62	: in std_logic := '0';
    EI63	: in std_logic := '0';
    EI64	: in std_logic := '0';
    EI65	: in std_logic := '0';
    EI66	: in std_logic := '0';
    EI67	: in std_logic := '0';
    EI68	: in std_logic := '0';
    EI69	: in std_logic := '0';
    EI70	: in std_logic := '0';
    EI71	: in std_logic := '0';
    EI72	: in std_logic := '0';
    EI73	: in std_logic := '0';
    EI74	: in std_logic := '0';
    EI75	: in std_logic := '0';
    EI76	: in std_logic := '0';
    EI77	: in std_logic := '0';
    EI78	: in std_logic := '0';
    EI79	: in std_logic := '0';
    EI80	: in std_logic := '0';
    EI81	: in std_logic := '0';
    EI82	: in std_logic := '0';
    EI83	: in std_logic := '0';
    EI84	: in std_logic := '0';
    EI85	: in std_logic := '0';
    EI86	: in std_logic := '0';
    EI87	: in std_logic := '0';
    EI88	: in std_logic := '0';
    EI89	: in std_logic := '0';
    EI90	: in std_logic := '0';
    EI91	: in std_logic := '0';
    EI92	: in std_logic := '0';
    EI93	: in std_logic := '0';
    EI94	: in std_logic := '0';
    EI95	: in std_logic := '0';
    EI96	: in std_logic := '0';
    EI97	: in std_logic := '0';
    EI98	: in std_logic := '0';
    EI99	: in std_logic := '0';
    EI100	: in std_logic := '0';
    EI101	: in std_logic := '0';
    EI102	: in std_logic := '0';
    EI103	: in std_logic := '0';
    EI104	: in std_logic := '0';
    EI105	: in std_logic := '0';
    EI106	: in std_logic := '0';
    EI107	: in std_logic := '0';
    EI108	: in std_logic := '0';
    EI109	: in std_logic := '0';
    EI110	: in std_logic := '0';
    EI111	: in std_logic := '0';
    EI112	: in std_logic := '0';
    EI113	: in std_logic := '0';
    EI114	: in std_logic := '0';
    EI115	: in std_logic := '0';
    EI116	: in std_logic := '0';
    EI117	: in std_logic := '0';
    EI118	: in std_logic := '0';
    EI119	: in std_logic := '0';
    EI120	: in std_logic := '0';
    EI121	: in std_logic := '0';
    EI122	: in std_logic := '0';
    EI123	: in std_logic := '0';
    EI124	: in std_logic := '0';
    EI125	: in std_logic := '0';
    EI126	: in std_logic := '0';
    EI127	: in std_logic := '0';
    EI128	: in std_logic := '0';
    EI129	: in std_logic := '0';
    EI130	: in std_logic := '0';
    EI131	: in std_logic := '0';
    EI132	: in std_logic := '0';
    EI133	: in std_logic := '0';
    EI134	: in std_logic := '0';
    EI135	: in std_logic := '0';
    EI136	: in std_logic := '0';
    EI137	: in std_logic := '0';
    EI138	: in std_logic := '0';
    EI139	: in std_logic := '0';
    EI140	: in std_logic := '0';
    EI141	: in std_logic := '0';
    EI142	: in std_logic := '0';
    EI143	: in std_logic := '0';
    EI144	: in std_logic := '0';
    EI145	: in std_logic := '0';
    EI146	: in std_logic := '0';
    EI147	: in std_logic := '0';
    EI148	: in std_logic := '0';
    EI149	: in std_logic := '0';
    EI150	: in std_logic := '0';
    EI151	: in std_logic := '0';
    EI152	: in std_logic := '0';
    EI153	: in std_logic := '0';
    EI154	: in std_logic := '0';
    EI155	: in std_logic := '0';
    EI156	: in std_logic := '0';
    EI157	: in std_logic := '0';
    EI158	: in std_logic := '0';
    EI159	: in std_logic := '0';
    EI160	: in std_logic := '0';
    EI161	: in std_logic := '0';
    EI162	: in std_logic := '0';
    EI163	: in std_logic := '0';
    EI164	: in std_logic := '0';
    EI165	: in std_logic := '0';
    EI166	: in std_logic := '0';
    EI167	: in std_logic := '0';
    EI168	: in std_logic := '0';
    EI169	: in std_logic := '0';
    EI170	: in std_logic := '0';
    EI171	: in std_logic := '0';
    EI172	: in std_logic := '0';
    EI173	: in std_logic := '0';
    EI174	: in std_logic := '0';
    EI175	: in std_logic := '0';
    EI176	: in std_logic := '0';
    EI177	: in std_logic := '0';
    EI178	: in std_logic := '0';
    EI179	: in std_logic := '0';
    EI180	: in std_logic := '0';
    EI181	: in std_logic := '0';
    EI182	: in std_logic := '0';
    EI183	: in std_logic := '0';
    EI184	: in std_logic := '0';
    EI185	: in std_logic := '0';
    EI186	: in std_logic := '0';
    EI187	: in std_logic := '0';
    EI188	: in std_logic := '0';
    EI189	: in std_logic := '0';
    EI190	: in std_logic := '0';
    EI191	: in std_logic := '0';
    EI192	: in std_logic := '0';
    EI_CK	: out std_logic := '0';
    EO_CK	: out std_logic := '0';
    EO1	: out std_logic := '0';
    EO2	: out std_logic := '0';
    EO3	: out std_logic := '0';
    EO4	: out std_logic := '0';
    EO5	: out std_logic := '0';
    EO6	: out std_logic := '0';
    EO7	: out std_logic := '0';
    EO8	: out std_logic := '0';
    EO9	: out std_logic := '0';
    EO10	: out std_logic := '0';
    EO11	: out std_logic := '0';
    EO12	: out std_logic := '0';
    EO13	: out std_logic := '0';
    EO14	: out std_logic := '0';
    EO15	: out std_logic := '0';
    EO16	: out std_logic := '0';
    EO17	: out std_logic := '0';
    EO18	: out std_logic := '0';
    EO19	: out std_logic := '0';
    EO20	: out std_logic := '0';
    EO21	: out std_logic := '0';
    EO22	: out std_logic := '0';
    EO23	: out std_logic := '0';
    EO24	: out std_logic := '0';
    EO25	: out std_logic := '0';
    EO26	: out std_logic := '0';
    EO27	: out std_logic := '0';
    EO28	: out std_logic := '0';
    EO29	: out std_logic := '0';
    EO30	: out std_logic := '0';
    EO31	: out std_logic := '0';
    EO32	: out std_logic := '0';
    EO33	: out std_logic := '0';
    EO34	: out std_logic := '0';
    EO35	: out std_logic := '0';
    EO36	: out std_logic := '0';
    EO37	: out std_logic := '0';
    EO38	: out std_logic := '0';
    EO39	: out std_logic := '0';
    EO40	: out std_logic := '0';
    EO41	: out std_logic := '0';
    EO42	: out std_logic := '0';
    EO43	: out std_logic := '0';
    EO44	: out std_logic := '0';
    EO45	: out std_logic := '0';
    EO46	: out std_logic := '0';
    EO47	: out std_logic := '0';
    EO48	: out std_logic := '0';
    EO49	: out std_logic := '0';
    EO50	: out std_logic := '0';
    EO51	: out std_logic := '0';
    EO52	: out std_logic := '0';
    EO53	: out std_logic := '0';
    EO54	: out std_logic := '0';
    EO55	: out std_logic := '0';
    EO56	: out std_logic := '0';
    EO57	: out std_logic := '0';
    EO58	: out std_logic := '0';
    EO59	: out std_logic := '0';
    EO60	: out std_logic := '0';
    EO61	: out std_logic := '0';
    EO62	: out std_logic := '0';
    EO63	: out std_logic := '0';
    EO64	: out std_logic := '0';
    EO65	: out std_logic := '0';
    EO66	: out std_logic := '0';
    EO67	: out std_logic := '0';
    EO68	: out std_logic := '0';
    EO69	: out std_logic := '0';
    EO70	: out std_logic := '0';
    EO71	: out std_logic := '0';
    EO72	: out std_logic := '0';
    EO73	: out std_logic := '0';
    EO74	: out std_logic := '0';
    EO75	: out std_logic := '0';
    EO76	: out std_logic := '0';
    EO77	: out std_logic := '0';
    EO78	: out std_logic := '0';
    EO79	: out std_logic := '0';
    EO80	: out std_logic := '0';
    EO81	: out std_logic := '0';
    EO82	: out std_logic := '0';
    EO83	: out std_logic := '0';
    EO84	: out std_logic := '0';
    EO85	: out std_logic := '0';
    EO86	: out std_logic := '0';
    EO87	: out std_logic := '0';
    EO88	: out std_logic := '0';
    EO89	: out std_logic := '0';
    EO90	: out std_logic := '0';
    EO91	: out std_logic := '0';
    EO92	: out std_logic := '0';
    EO93	: out std_logic := '0';
    EO94	: out std_logic := '0';
    EO95	: out std_logic := '0';
    EO96	: out std_logic := '0';
    EO97	: out std_logic := '0';
    EO98	: out std_logic := '0';
    EO99	: out std_logic := '0';
    EO100	: out std_logic := '0';
    EO101	: out std_logic := '0';
    EO102	: out std_logic := '0';
    EO103	: out std_logic := '0';
    EO104	: out std_logic := '0';
    EO105	: out std_logic := '0';
    EO106	: out std_logic := '0';
    EO107	: out std_logic := '0';
    EO108	: out std_logic := '0';
    EO109	: out std_logic := '0';
    EO110	: out std_logic := '0';
    EO111	: out std_logic := '0';
    EO112	: out std_logic := '0';
    EO113	: out std_logic := '0';
    EO114	: out std_logic := '0';
    EO115	: out std_logic := '0';
    EO116	: out std_logic := '0';
    EO117	: out std_logic := '0';
    EO118	: out std_logic := '0';
    EO119	: out std_logic := '0';
    EO120	: out std_logic := '0';
    EO121	: out std_logic := '0';
    EO122	: out std_logic := '0';
    EO123	: out std_logic := '0';
    EO124	: out std_logic := '0';
    EO125	: out std_logic := '0';
    EO126	: out std_logic := '0';
    EO127	: out std_logic := '0';
    EO128	: out std_logic := '0';
    EO129	: out std_logic := '0';
    EO130	: out std_logic := '0';
    EO131	: out std_logic := '0';
    EO132	: out std_logic := '0';
    EO133	: out std_logic := '0';
    EO134	: out std_logic := '0';
    EO135	: out std_logic := '0';
    EO136	: out std_logic := '0';
    EO137	: out std_logic := '0';
    EO138	: out std_logic := '0';
    EO139	: out std_logic := '0';
    EO140	: out std_logic := '0';
    EO141	: out std_logic := '0';
    EO142	: out std_logic := '0';
    EO143	: out std_logic := '0';
    EO144	: out std_logic := '0';
    EO145	: out std_logic := '0';
    EO146	: out std_logic := '0';
    EO147	: out std_logic := '0';
    EO148	: out std_logic := '0';
    EO149	: out std_logic := '0';
    EO150	: out std_logic := '0';
    EO151	: out std_logic := '0';
    EO152	: out std_logic := '0';
    EO153	: out std_logic := '0';
    EO154	: out std_logic := '0';
    EO155	: out std_logic := '0';
    EO156	: out std_logic := '0';
    EO157	: out std_logic := '0';
    EO158	: out std_logic := '0';
    EO159	: out std_logic := '0';
    EO160	: out std_logic := '0';
    EO161	: out std_logic := '0';
    EO162	: out std_logic := '0';
    EO163	: out std_logic := '0';
    EO164	: out std_logic := '0';
    EO165	: out std_logic := '0';
    EO166	: out std_logic := '0';
    EO167	: out std_logic := '0';
    EO168	: out std_logic := '0';
    EO169	: out std_logic := '0';
    EO170	: out std_logic := '0';
    EO171	: out std_logic := '0';
    EO172	: out std_logic := '0';
    EO173	: out std_logic := '0';
    EO174	: out std_logic := '0';
    EO175	: out std_logic := '0';
    EO176	: out std_logic := '0';
    EO177	: out std_logic := '0';
    EO178	: out std_logic := '0';
    EO179	: out std_logic := '0';
    EO180	: out std_logic := '0';
    EO181	: out std_logic := '0';
    EO182	: out std_logic := '0';
    EO183	: out std_logic := '0';
    EO184	: out std_logic := '0';
    EO185	: out std_logic := '0';
    EO186	: out std_logic := '0';
    EO187	: out std_logic := '0';
    EO188	: out std_logic := '0';
    EO189	: out std_logic := '0';
    EO190	: out std_logic := '0';
    EO191	: out std_logic := '0';
    EO192	: out std_logic := '0';
    FI1	: in std_logic := '0';
    FI2	: in std_logic := '0';
    FI3	: in std_logic := '0';
    FI4	: in std_logic := '0';
    FI5	: in std_logic := '0';
    FI6	: in std_logic := '0';
    FI7	: in std_logic := '0';
    FI8	: in std_logic := '0';
    FI9	: in std_logic := '0';
    FI10	: in std_logic := '0';
    FI11	: in std_logic := '0';
    FI12	: in std_logic := '0';
    FI13	: in std_logic := '0';
    FI14	: in std_logic := '0';
    FI15	: in std_logic := '0';
    FI16	: in std_logic := '0';
    FI17	: in std_logic := '0';
    FI18	: in std_logic := '0';
    FI19	: in std_logic := '0';
    FI20	: in std_logic := '0';
    FI21	: in std_logic := '0';
    FI22	: in std_logic := '0';
    FI23	: in std_logic := '0';
    FI24	: in std_logic := '0';
    FI25	: in std_logic := '0';
    FI26	: in std_logic := '0';
    FI27	: in std_logic := '0';
    FI28	: in std_logic := '0';
    FI29	: in std_logic := '0';
    FI30	: in std_logic := '0';
    FI31	: in std_logic := '0';
    FI32	: in std_logic := '0';
    FI33	: in std_logic := '0';
    FI34	: in std_logic := '0';
    FI35	: in std_logic := '0';
    FI36	: in std_logic := '0';
    FI37	: in std_logic := '0';
    FI38	: in std_logic := '0';
    FI39	: in std_logic := '0';
    FI40	: in std_logic := '0';
    FI41	: in std_logic := '0';
    FI42	: in std_logic := '0';
    FI43	: in std_logic := '0';
    FI44	: in std_logic := '0';
    FI45	: in std_logic := '0';
    FI46	: in std_logic := '0';
    FI47	: in std_logic := '0';
    FI48	: in std_logic := '0';
    FI49	: in std_logic := '0';
    FI50	: in std_logic := '0';
    FI51	: in std_logic := '0';
    FI52	: in std_logic := '0';
    FI53	: in std_logic := '0';
    FI54	: in std_logic := '0';
    FI55	: in std_logic := '0';
    FI56	: in std_logic := '0';
    FI57	: in std_logic := '0';
    FI58	: in std_logic := '0';
    FI59	: in std_logic := '0';
    FI60	: in std_logic := '0';
    FI61	: in std_logic := '0';
    FI62	: in std_logic := '0';
    FI63	: in std_logic := '0';
    FI64	: in std_logic := '0';
    FI65	: in std_logic := '0';
    FI66	: in std_logic := '0';
    FI67	: in std_logic := '0';
    FI68	: in std_logic := '0';
    FI69	: in std_logic := '0';
    FI70	: in std_logic := '0';
    FI71	: in std_logic := '0';
    FI72	: in std_logic := '0';
    FI73	: in std_logic := '0';
    FI74	: in std_logic := '0';
    FI75	: in std_logic := '0';
    FI76	: in std_logic := '0';
    FI77	: in std_logic := '0';
    FI78	: in std_logic := '0';
    FI79	: in std_logic := '0';
    FI80	: in std_logic := '0';
    FI81	: in std_logic := '0';
    FI82	: in std_logic := '0';
    FI83	: in std_logic := '0';
    FI84	: in std_logic := '0';
    FI85	: in std_logic := '0';
    FI86	: in std_logic := '0';
    FI87	: in std_logic := '0';
    FI88	: in std_logic := '0';
    FI89	: in std_logic := '0';
    FI90	: in std_logic := '0';
    FI91	: in std_logic := '0';
    FI92	: in std_logic := '0';
    FI93	: in std_logic := '0';
    FI94	: in std_logic := '0';
    FI95	: in std_logic := '0';
    FI96	: in std_logic := '0';
    FI97	: in std_logic := '0';
    FI98	: in std_logic := '0';
    FI99	: in std_logic := '0';
    FI100	: in std_logic := '0';
    FI101	: in std_logic := '0';
    FI102	: in std_logic := '0';
    FI103	: in std_logic := '0';
    FI104	: in std_logic := '0';
    FI105	: in std_logic := '0';
    FI106	: in std_logic := '0';
    FI107	: in std_logic := '0';
    FI108	: in std_logic := '0';
    FI109	: in std_logic := '0';
    FI110	: in std_logic := '0';
    FI111	: in std_logic := '0';
    FI112	: in std_logic := '0';
    FI113	: in std_logic := '0';
    FI114	: in std_logic := '0';
    FI115	: in std_logic := '0';
    FI116	: in std_logic := '0';
    FI117	: in std_logic := '0';
    FI118	: in std_logic := '0';
    FI119	: in std_logic := '0';
    FI120	: in std_logic := '0';
    FI121	: in std_logic := '0';
    FI122	: in std_logic := '0';
    FI123	: in std_logic := '0';
    FI124	: in std_logic := '0';
    FI125	: in std_logic := '0';
    FI126	: in std_logic := '0';
    FI127	: in std_logic := '0';
    FI128	: in std_logic := '0';
    FI129	: in std_logic := '0';
    FI130	: in std_logic := '0';
    FI131	: in std_logic := '0';
    FI132	: in std_logic := '0';
    FI133	: in std_logic := '0';
    FI134	: in std_logic := '0';
    FI135	: in std_logic := '0';
    FI136	: in std_logic := '0';
    FI137	: in std_logic := '0';
    FI138	: in std_logic := '0';
    FI139	: in std_logic := '0';
    FI140	: in std_logic := '0';
    FI141	: in std_logic := '0';
    FI142	: in std_logic := '0';
    FI143	: in std_logic := '0';
    FI144	: in std_logic := '0';
    FI145	: in std_logic := '0';
    FI146	: in std_logic := '0';
    FI147	: in std_logic := '0';
    FI148	: in std_logic := '0';
    FI149	: in std_logic := '0';
    FI150	: in std_logic := '0';
    FI151	: in std_logic := '0';
    FI152	: in std_logic := '0';
    FI153	: in std_logic := '0';
    FI154	: in std_logic := '0';
    FI155	: in std_logic := '0';
    FI156	: in std_logic := '0';
    FI157	: in std_logic := '0';
    FI158	: in std_logic := '0';
    FI159	: in std_logic := '0';
    FI160	: in std_logic := '0';
    FI161	: in std_logic := '0';
    FI162	: in std_logic := '0';
    FI163	: in std_logic := '0';
    FI164	: in std_logic := '0';
    FI165	: in std_logic := '0';
    FI166	: in std_logic := '0';
    FI167	: in std_logic := '0';
    FI168	: in std_logic := '0';
    FI169	: in std_logic := '0';
    FI170	: in std_logic := '0';
    FI171	: in std_logic := '0';
    FI172	: in std_logic := '0';
    FI173	: in std_logic := '0';
    FI174	: in std_logic := '0';
    FI175	: in std_logic := '0';
    FI176	: in std_logic := '0';
    FI177	: in std_logic := '0';
    FI178	: in std_logic := '0';
    FI179	: in std_logic := '0';
    FI180	: in std_logic := '0';
    FI181	: in std_logic := '0';
    FI182	: in std_logic := '0';
    FI183	: in std_logic := '0';
    FI184	: in std_logic := '0';
    FI185	: in std_logic := '0';
    FI186	: in std_logic := '0';
    FI187	: in std_logic := '0';
    FI188	: in std_logic := '0';
    FI189	: in std_logic := '0';
    FI190	: in std_logic := '0';
    FI191	: in std_logic := '0';
    FI192	: in std_logic := '0';
    FO1	: out std_logic := '0';
    FO2	: out std_logic := '0';
    FO3	: out std_logic := '0';
    FO4	: out std_logic := '0';
    FO5	: out std_logic := '0';
    FO6	: out std_logic := '0';
    FO7	: out std_logic := '0';
    FO8	: out std_logic := '0';
    FO9	: out std_logic := '0';
    FO10	: out std_logic := '0';
    FO11	: out std_logic := '0';
    FO12	: out std_logic := '0';
    FO13	: out std_logic := '0';
    FO14	: out std_logic := '0';
    FO15	: out std_logic := '0';
    FO16	: out std_logic := '0';
    FO17	: out std_logic := '0';
    FO18	: out std_logic := '0';
    FO19	: out std_logic := '0';
    FO20	: out std_logic := '0';
    FO21	: out std_logic := '0';
    FO22	: out std_logic := '0';
    FO23	: out std_logic := '0';
    FO24	: out std_logic := '0';
    FO25	: out std_logic := '0';
    FO26	: out std_logic := '0';
    FO27	: out std_logic := '0';
    FO28	: out std_logic := '0';
    FO29	: out std_logic := '0';
    FO30	: out std_logic := '0';
    FO31	: out std_logic := '0';
    FO32	: out std_logic := '0';
    FO33	: out std_logic := '0';
    FO34	: out std_logic := '0';
    FO35	: out std_logic := '0';
    FO36	: out std_logic := '0';
    FO37	: out std_logic := '0';
    FO38	: out std_logic := '0';
    FO39	: out std_logic := '0';
    FO40	: out std_logic := '0';
    FO41	: out std_logic := '0';
    FO42	: out std_logic := '0';
    FO43	: out std_logic := '0';
    FO44	: out std_logic := '0';
    FO45	: out std_logic := '0';
    FO46	: out std_logic := '0';
    FO47	: out std_logic := '0';
    FO48	: out std_logic := '0';
    FO49	: out std_logic := '0';
    FO50	: out std_logic := '0';
    FO51	: out std_logic := '0';
    FO52	: out std_logic := '0';
    FO53	: out std_logic := '0';
    FO54	: out std_logic := '0';
    FO55	: out std_logic := '0';
    FO56	: out std_logic := '0';
    FO57	: out std_logic := '0';
    FO58	: out std_logic := '0';
    FO59	: out std_logic := '0';
    FO60	: out std_logic := '0';
    FO61	: out std_logic := '0';
    FO62	: out std_logic := '0';
    FO63	: out std_logic := '0';
    FO64	: out std_logic := '0';
    FO65	: out std_logic := '0';
    FO66	: out std_logic := '0';
    FO67	: out std_logic := '0';
    FO68	: out std_logic := '0';
    FO69	: out std_logic := '0';
    FO70	: out std_logic := '0';
    FO71	: out std_logic := '0';
    FO72	: out std_logic := '0';
    FO73	: out std_logic := '0';
    FO74	: out std_logic := '0';
    FO75	: out std_logic := '0';
    FO76	: out std_logic := '0';
    FO77	: out std_logic := '0';
    FO78	: out std_logic := '0';
    FO79	: out std_logic := '0';
    FO80	: out std_logic := '0';
    FO81	: out std_logic := '0';
    FO82	: out std_logic := '0';
    FO83	: out std_logic := '0';
    FO84	: out std_logic := '0';
    FO85	: out std_logic := '0';
    FO86	: out std_logic := '0';
    FO87	: out std_logic := '0';
    FO88	: out std_logic := '0';
    FO89	: out std_logic := '0';
    FO90	: out std_logic := '0';
    FO91	: out std_logic := '0';
    FO92	: out std_logic := '0';
    FO93	: out std_logic := '0';
    FO94	: out std_logic := '0';
    FO95	: out std_logic := '0';
    FO96	: out std_logic := '0';
    FO97	: out std_logic := '0';
    FO98	: out std_logic := '0';
    FO99	: out std_logic := '0';
    FO100	: out std_logic := '0';
    FO101	: out std_logic := '0';
    FO102	: out std_logic := '0';
    FO103	: out std_logic := '0';
    FO104	: out std_logic := '0';
    FO105	: out std_logic := '0';
    FO106	: out std_logic := '0';
    FO107	: out std_logic := '0';
    FO108	: out std_logic := '0';
    FO109	: out std_logic := '0';
    FO110	: out std_logic := '0';
    FO111	: out std_logic := '0';
    FO112	: out std_logic := '0';
    FO113	: out std_logic := '0';
    FO114	: out std_logic := '0';
    FO115	: out std_logic := '0';
    FO116	: out std_logic := '0';
    FO117	: out std_logic := '0';
    FO118	: out std_logic := '0';
    FO119	: out std_logic := '0';
    FO120	: out std_logic := '0';
    FO121	: out std_logic := '0';
    FO122	: out std_logic := '0';
    FO123	: out std_logic := '0';
    FO124	: out std_logic := '0';
    FO125	: out std_logic := '0';
    FO126	: out std_logic := '0';
    FO127	: out std_logic := '0';
    FO128	: out std_logic := '0';
    FO129	: out std_logic := '0';
    FO130	: out std_logic := '0';
    FO131	: out std_logic := '0';
    FO132	: out std_logic := '0';
    FO133	: out std_logic := '0';
    FO134	: out std_logic := '0';
    FO135	: out std_logic := '0';
    FO136	: out std_logic := '0';
    FO137	: out std_logic := '0';
    FO138	: out std_logic := '0';
    FO139	: out std_logic := '0';
    FO140	: out std_logic := '0';
    FO141	: out std_logic := '0';
    FO142	: out std_logic := '0';
    FO143	: out std_logic := '0';
    FO144	: out std_logic := '0';
    FO145	: out std_logic := '0';
    FO146	: out std_logic := '0';
    FO147	: out std_logic := '0';
    FO148	: out std_logic := '0';
    FO149	: out std_logic := '0';
    FO150	: out std_logic := '0';
    FO151	: out std_logic := '0';
    FO152	: out std_logic := '0';
    FO153	: out std_logic := '0';
    FO154	: out std_logic := '0';
    FO155	: out std_logic := '0';
    FO156	: out std_logic := '0';
    FO157	: out std_logic := '0';
    FO158	: out std_logic := '0';
    FO159	: out std_logic := '0';
    FO160	: out std_logic := '0';
    FO161	: out std_logic := '0';
    FO162	: out std_logic := '0';
    FO163	: out std_logic := '0';
    FO164	: out std_logic := '0';
    FO165	: out std_logic := '0';
    FO166	: out std_logic := '0';
    FO167	: out std_logic := '0';
    FO168	: out std_logic := '0';
    FO169	: out std_logic := '0';
    FO170	: out std_logic := '0';
    FO171	: out std_logic := '0';
    FO172	: out std_logic := '0';
    FO173	: out std_logic := '0';
    FO174	: out std_logic := '0';
    FO175	: out std_logic := '0';
    FO176	: out std_logic := '0';
    FO177	: out std_logic := '0';
    FO178	: out std_logic := '0';
    FO179	: out std_logic := '0';
    FO180	: out std_logic := '0';
    FO181	: out std_logic := '0';
    FO182	: out std_logic := '0';
    FO183	: out std_logic := '0';
    FO184	: out std_logic := '0';
    FO185	: out std_logic := '0';
    FO186	: out std_logic := '0';
    FO187	: out std_logic := '0';
    FO188	: out std_logic := '0';
    FO189	: out std_logic := '0';
    FO190	: out std_logic := '0';
    FO191	: out std_logic := '0';
    FO192	: out std_logic := '0'
);
end component NX_RB;

component NX_RB_WRAP is
generic (
    -- input : EI to FO
    inputClk      : bit_vector( 1 downto 0) := B"00"; -- 00 = CK[0], 01 = CK[1], 10 = CK[2] and 11 = CK[3]
    inputBypass   : bit_vector(23 downto 0) := B"000000000000000000000000"; -- 1 bypass active, LSB is bypass registers 0 to 7 ... MSB is bypass registers 183 to 191
    -- output : FI to EO
    inputContext  : string := ""; -- input context intialization
    outputClk     : bit_vector( 1 downto 0) := B"00"; -- 00 = CK[0], 01 = CK[1], 10 = CK[2] and 11 = CK[3]
    outputBypass  : bit_vector(23 downto 0) := B"000000000000000000000000";  -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    outputContext : string := "" -- output context intialization
);
port (
    CK	: in std_logic_vector(  3 downto 0) := (others => '0');
    EI_CK	: out std_logic := '0';
    EO_CK	: out std_logic := '0';
    EI	: in std_logic_vector(191 downto 0) := (others => '0');
    EO	: out std_logic_vector(191 downto 0) := (others => '0');
    FI	: in std_logic_vector(191 downto 0) := (others => '0');
    FO	: out std_logic_vector(191 downto 0) := (others => '0')
);
end component NX_RB_WRAP;

component NX_RFB_L is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    I5	: in std_logic := '0';
    I6	: in std_logic := '0';
    I7	: in std_logic := '0';
    I8	: in std_logic := '0';
    I9	: in std_logic := '0';
    I10	: in std_logic := '0';
    I11	: in std_logic := '0';
    I12	: in std_logic := '0';
    I13	: in std_logic := '0';
    I14	: in std_logic := '0';
    I15	: in std_logic := '0';
    I16	: in std_logic := '0';
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0';
    O1	: out std_logic := '0';
    O2	: out std_logic := '0';
    O3	: out std_logic := '0';
    O4	: out std_logic := '0';
    O5	: out std_logic := '0';
    O6	: out std_logic := '0';
    O7	: out std_logic := '0';
    O8	: out std_logic := '0';
    O9	: out std_logic := '0';
    O10	: out std_logic := '0';
    O11	: out std_logic := '0';
    O12	: out std_logic := '0';
    O13	: out std_logic := '0';
    O14	: out std_logic := '0';
    O15	: out std_logic := '0';
    O16	: out std_logic := '0';
    RA1	: in std_logic := '0';
    RA2	: in std_logic := '0';
    RA3	: in std_logic := '0';
    RA4	: in std_logic := '0';
    RA5	: in std_logic := '0';
    RA6	: in std_logic := '0';
    RE	: in std_logic := '0';
    WA1	: in std_logic := '0';
    WA2	: in std_logic := '0';
    WA3	: in std_logic := '0';
    WA4	: in std_logic := '0';
    WA5	: in std_logic := '0';
    WA6	: in std_logic := '0';
    WE	: in std_logic := '0';
    XRCK	: out std_logic := '0';
    XRO1	: out std_logic := '0';
    XRO2	: out std_logic := '0';
    XRO3	: out std_logic := '0';
    XRO4	: out std_logic := '0';
    XRO5	: out std_logic := '0';
    XRO6	: out std_logic := '0';
    XWCK	: out std_logic := '0';
    XWO1	: out std_logic := '0';
    XWO2	: out std_logic := '0';
    XWO3	: out std_logic := '0';
    XWO4	: out std_logic := '0';
    XWO5	: out std_logic := '0';
    XWO6	: out std_logic := '0'
);
end component NX_RFB_L;

component NX_RFB_L_WRAP is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(15 downto 0) := (others => '0');
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0';
    O	: out std_logic_vector(15 downto 0) := (others => '0');
    RA	: in std_logic_vector(5 downto 0) := (others => '0');
    RE	: in std_logic := '0';
    WA	: in std_logic_vector(5 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    XRCK	: out std_logic := '0';
    XRO	: out std_logic_vector(5 downto 0) := (others => '0');
    XWCK	: out std_logic := '0';
    XWO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_RFB_L_WRAP;

component NX_RFB_M is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    I5	: in std_logic := '0';
    I6	: in std_logic := '0';
    I7	: in std_logic := '0';
    I8	: in std_logic := '0';
    I9	: in std_logic := '0';
    I10	: in std_logic := '0';
    I11	: in std_logic := '0';
    I12	: in std_logic := '0';
    I13	: in std_logic := '0';
    I14	: in std_logic := '0';
    I15	: in std_logic := '0';
    I16	: in std_logic := '0';
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0';
    O1	: out std_logic := '0';
    O2	: out std_logic := '0';
    O3	: out std_logic := '0';
    O4	: out std_logic := '0';
    O5	: out std_logic := '0';
    O6	: out std_logic := '0';
    O7	: out std_logic := '0';
    O8	: out std_logic := '0';
    O9	: out std_logic := '0';
    O10	: out std_logic := '0';
    O11	: out std_logic := '0';
    O12	: out std_logic := '0';
    O13	: out std_logic := '0';
    O14	: out std_logic := '0';
    O15	: out std_logic := '0';
    O16	: out std_logic := '0';
    RA1	: in std_logic := '0';
    RA2	: in std_logic := '0';
    RA3	: in std_logic := '0';
    RA4	: in std_logic := '0';
    RA5	: in std_logic := '0';
    RA6	: in std_logic := '0';
    RE	: in std_logic := '0';
    WA1	: in std_logic := '0';
    WA2	: in std_logic := '0';
    WA3	: in std_logic := '0';
    WA4	: in std_logic := '0';
    WA5	: in std_logic := '0';
    WA6	: in std_logic := '0';
    WE	: in std_logic := '0'
);
end component NX_RFB_M;

component NX_RFB_WRAP is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(15 downto 0) := (others => '0');
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0';
    O	: out std_logic_vector(15 downto 0) := (others => '0');
    RA	: in std_logic_vector(5 downto 0) := (others => '0');
    RE	: in std_logic := '0';
    WA	: in std_logic_vector(5 downto 0) := (others => '0');
    WE	: in std_logic := '0'
);
end component NX_RFB_WRAP;

component NX_CKS is
port (
    CKI	: in std_logic := '0';
    CMD	: in std_logic := '0';
    CKO	: out std_logic := '0'
);
end component NX_CKS;

component NX_RFB is
generic (
    rck_edge  : bit := '0';   -- 0: read  clock rising edge - 1: read  clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK	: in std_logic := '0';
    WCK	: in std_logic := '0';
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    I5	: in std_logic := '0';
    I6	: in std_logic := '0';
    I7	: in std_logic := '0';
    I8	: in std_logic := '0';
    I9	: in std_logic := '0';
    I10	: in std_logic := '0';
    I11	: in std_logic := '0';
    I12	: in std_logic := '0';
    I13	: in std_logic := '0';
    I14	: in std_logic := '0';
    I15	: in std_logic := '0';
    I16	: in std_logic := '0';
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0';
    O1	: out std_logic := '0';
    O2	: out std_logic := '0';
    O3	: out std_logic := '0';
    O4	: out std_logic := '0';
    O5	: out std_logic := '0';
    O6	: out std_logic := '0';
    O7	: out std_logic := '0';
    O8	: out std_logic := '0';
    O9	: out std_logic := '0';
    O10	: out std_logic := '0';
    O11	: out std_logic := '0';
    O12	: out std_logic := '0';
    O13	: out std_logic := '0';
    O14	: out std_logic := '0';
    O15	: out std_logic := '0';
    O16	: out std_logic := '0';
    RA1	: in std_logic := '0';
    RA2	: in std_logic := '0';
    RA3	: in std_logic := '0';
    RA4	: in std_logic := '0';
    RA5	: in std_logic := '0';
    RA6	: in std_logic := '0';
    RE	: in std_logic := '0';
    WA1	: in std_logic := '0';
    WA2	: in std_logic := '0';
    WA3	: in std_logic := '0';
    WA4	: in std_logic := '0';
    WA5	: in std_logic := '0';
    WA6	: in std_logic := '0';
    WE	: in std_logic := '0'
);
end component NX_RFB;

component NX_CDC_U_2DFF is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_adest_arst : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    ADRSTI	: in std_logic := '0';
    ADRSTO	: out std_logic := '0';
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BDRSTI	: in std_logic := '0';
    BDRSTO	: out std_logic := '0';
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_CDC_U_2DFF;

component NX_CDC_U_3DFF is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    ASRSTI	: in std_logic := '0';
    ADRSTI	: in std_logic := '0';
    ASRSTO	: out std_logic := '0';
    ADRSTO	: out std_logic := '0';
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BSRSTI	: in std_logic := '0';
    BDRSTI	: in std_logic := '0';
    BSRSTO	: out std_logic := '0';
    BDRSTO	: out std_logic := '0';
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_CDC_U_3DFF;

component NX_CDC_U_FULL is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    ASRSTI	: in std_logic := '0';
    ADRSTI	: in std_logic := '0';
    ASRSTO	: out std_logic := '0';
    ADRSTO	: out std_logic := '0';
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BSRSTI	: in std_logic := '0';
    BDRSTI	: in std_logic := '0';
    BSRSTO	: out std_logic := '0';
    BDRSTO	: out std_logic := '0';
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_CDC_U_FULL;

component NX_CDC_U_BIN2GRAY is
port (
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_CDC_U_BIN2GRAY;

component NX_CDC_U_GRAY2BIN is
port (
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_CDC_U_GRAY2BIN;

component NX_XCDC_U is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    ASRSTI	: in std_logic := '0';
    ADRSTI	: in std_logic := '0';
    ASRSTO	: out std_logic := '0';
    ADRSTO	: out std_logic := '0';
    AI	: in std_logic_vector(5 downto 0) := (others => '0');
    AO	: out std_logic_vector(5 downto 0) := (others => '0');
    BSRSTI	: in std_logic := '0';
    BDRSTI	: in std_logic := '0';
    BSRSTO	: out std_logic := '0';
    BDRSTO	: out std_logic := '0';
    BI	: in std_logic_vector(5 downto 0) := (others => '0');
    BO	: out std_logic_vector(5 downto 0) := (others => '0');
    CSRSTI	: in std_logic := '0';
    CDRSTI	: in std_logic := '0';
    CSRSTO	: out std_logic := '0';
    CDRSTO	: out std_logic := '0';
    CI	: in std_logic_vector(5 downto 0) := (others => '0');
    CO	: out std_logic_vector(5 downto 0) := (others => '0');
    DSRSTI	: in std_logic := '0';
    DDRSTI	: in std_logic := '0';
    DSRSTO	: out std_logic := '0';
    DDRSTO	: out std_logic := '0';
    DI	: in std_logic_vector(5 downto 0) := (others => '0');
    DO	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_XCDC_U;

component NX_CDC_U is
generic (
    mode           : integer := 0; -- 0: 2DFF     
                                   -- 1: 3DFF     
                                   -- 2: bin2gray + 3DFF + gray2bin
                                   -- 3: bin2gray 
                                   -- 4: gray2bin 
                                   -- 5: XCDC
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1	: in std_logic := '0';
    CK2	: in std_logic := '0';
    ASRSTI	: in std_logic := '0';
    ADRSTI	: in std_logic := '0';
    ASRSTO	: out std_logic := '0';
    ADRSTO	: out std_logic := '0';
    AI1	: in std_logic := '0';
    AI2	: in std_logic := '0';
    AI3	: in std_logic := '0';
    AI4	: in std_logic := '0';
    AI5	: in std_logic := '0';
    AI6	: in std_logic := '0';
    AO1	: out std_logic := '0';
    AO2	: out std_logic := '0';
    AO3	: out std_logic := '0';
    AO4	: out std_logic := '0';
    AO5	: out std_logic := '0';
    AO6	: out std_logic := '0';
    BSRSTI	: in std_logic := '0';
    BDRSTI	: in std_logic := '0';
    BSRSTO	: out std_logic := '0';
    BDRSTO	: out std_logic := '0';
    BI1	: in std_logic := '0';
    BI2	: in std_logic := '0';
    BI3	: in std_logic := '0';
    BI4	: in std_logic := '0';
    BI5	: in std_logic := '0';
    BI6	: in std_logic := '0';
    BO1	: out std_logic := '0';
    BO2	: out std_logic := '0';
    BO3	: out std_logic := '0';
    BO4	: out std_logic := '0';
    BO5	: out std_logic := '0';
    BO6	: out std_logic := '0';
    CSRSTI	: in std_logic := '0';
    CDRSTI	: in std_logic := '0';
    CSRSTO	: out std_logic := '0';
    CDRSTO	: out std_logic := '0';
    CI1	: in std_logic := '0';
    CI2	: in std_logic := '0';
    CI3	: in std_logic := '0';
    CI4	: in std_logic := '0';
    CI5	: in std_logic := '0';
    CI6	: in std_logic := '0';
    CO1	: out std_logic := '0';
    CO2	: out std_logic := '0';
    CO3	: out std_logic := '0';
    CO4	: out std_logic := '0';
    CO5	: out std_logic := '0';
    CO6	: out std_logic := '0';
    DSRSTI	: in std_logic := '0';
    DDRSTI	: in std_logic := '0';
    DSRSTO	: out std_logic := '0';
    DDRSTO	: out std_logic := '0';
    DI1	: in std_logic := '0';
    DI2	: in std_logic := '0';
    DI3	: in std_logic := '0';
    DI4	: in std_logic := '0';
    DI5	: in std_logic := '0';
    DI6	: in std_logic := '0';
    DO1	: out std_logic := '0';
    DO2	: out std_logic := '0';
    DO3	: out std_logic := '0';
    DO4	: out std_logic := '0';
    DO5	: out std_logic := '0';
    DO6	: out std_logic := '0'
);
end component NX_CDC_U;

component NX_RFB_U_WRAP is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    O	: out std_logic_vector(17 downto 0) := (others => '0');
    RA	: in std_logic_vector(4 downto 0) := (others => '0');
    WA	: in std_logic_vector(4 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_RFB_U_WRAP;

component NX_RFBSP_U_WRAP is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    O	: out std_logic_vector(17 downto 0) := (others => '0');
    WA	: in std_logic_vector(4 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_RFBSP_U_WRAP;

component NX_RFB_U is
generic (
    mode     : integer := 0; -- 0: DPREG - 1: SPREG - 2: XRF_64x18 - 3: XRF_32x36 - 4: XRF_2R_1W
    wck_edge : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    I5	: in std_logic := '0';
    I6	: in std_logic := '0';
    I7	: in std_logic := '0';
    I8	: in std_logic := '0';
    I9	: in std_logic := '0';
    I10	: in std_logic := '0';
    I11	: in std_logic := '0';
    I12	: in std_logic := '0';
    I13	: in std_logic := '0';
    I14	: in std_logic := '0';
    I15	: in std_logic := '0';
    I16	: in std_logic := '0';
    I17	: in std_logic := '0';
    I18	: in std_logic := '0';
    I19	: in std_logic := '0';
    I20	: in std_logic := '0';
    I21	: in std_logic := '0';
    I22	: in std_logic := '0';
    I23	: in std_logic := '0';
    I24	: in std_logic := '0';
    I25	: in std_logic := '0';
    I26	: in std_logic := '0';
    I27	: in std_logic := '0';
    I28	: in std_logic := '0';
    I29	: in std_logic := '0';
    I30	: in std_logic := '0';
    I31	: in std_logic := '0';
    I32	: in std_logic := '0';
    I33	: in std_logic := '0';
    I34	: in std_logic := '0';
    I35	: in std_logic := '0';
    I36	: in std_logic := '0';
    O1	: out std_logic := '0';
    O2	: out std_logic := '0';
    O3	: out std_logic := '0';
    O4	: out std_logic := '0';
    O5	: out std_logic := '0';
    O6	: out std_logic := '0';
    O7	: out std_logic := '0';
    O8	: out std_logic := '0';
    O9	: out std_logic := '0';
    O10	: out std_logic := '0';
    O11	: out std_logic := '0';
    O12	: out std_logic := '0';
    O13	: out std_logic := '0';
    O14	: out std_logic := '0';
    O15	: out std_logic := '0';
    O16	: out std_logic := '0';
    O17	: out std_logic := '0';
    O18	: out std_logic := '0';
    O19	: out std_logic := '0';
    O20	: out std_logic := '0';
    O21	: out std_logic := '0';
    O22	: out std_logic := '0';
    O23	: out std_logic := '0';
    O24	: out std_logic := '0';
    O25	: out std_logic := '0';
    O26	: out std_logic := '0';
    O27	: out std_logic := '0';
    O28	: out std_logic := '0';
    O29	: out std_logic := '0';
    O30	: out std_logic := '0';
    O31	: out std_logic := '0';
    O32	: out std_logic := '0';
    O33	: out std_logic := '0';
    O34	: out std_logic := '0';
    O35	: out std_logic := '0';
    O36	: out std_logic := '0';
    RA1	: in std_logic := '0';
    RA2	: in std_logic := '0';
    RA3	: in std_logic := '0';
    RA4	: in std_logic := '0';
    RA5	: in std_logic := '0';
    RA6	: in std_logic := '0';
    RA7	: in std_logic := '0';
    RA8	: in std_logic := '0';
    RA9	: in std_logic := '0';
    RA10	: in std_logic := '0';
    WA1	: in std_logic := '0';
    WA2	: in std_logic := '0';
    WA3	: in std_logic := '0';
    WA4	: in std_logic := '0';
    WA5	: in std_logic := '0';
    WA6	: in std_logic := '0';
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_RFB_U;

component NX_XRFB_64x18 is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    O	: out std_logic_vector(17 downto 0) := (others => '0');
    RA	: in std_logic_vector(5 downto 0) := (others => '0');
    WA	: in std_logic_vector(5 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_XRFB_64x18;

component NX_XRFB_32x36 is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(35 downto 0) := (others => '0');
    O	: out std_logic_vector(35 downto 0) := (others => '0');
    RA	: in std_logic_vector(4 downto 0) := (others => '0');
    WA	: in std_logic_vector(4 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_XRFB_32x36;

component NX_XRFB_2R_1W is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK	: in std_logic := '0';
    I	: in std_logic_vector(17 downto 0) := (others => '0');
    AO	: out std_logic_vector(17 downto 0) := (others => '0');
    BO	: out std_logic_vector(17 downto 0) := (others => '0');
    ARA	: in std_logic_vector(4 downto 0) := (others => '0');
    BRA	: in std_logic_vector(4 downto 0) := (others => '0');
    WA	: in std_logic_vector(4 downto 0) := (others => '0');
    WE	: in std_logic := '0';
    WEA	: in std_logic := '0'
);
end component NX_XRFB_2R_1W;

component NX_SER is
generic (
    data_size            : integer range 2 to 10 := 5;	-- Number of serialization factor
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0") or differential ("1")
    slewRate             : string := "";		-- Slow, Medium or Fast
    outputDelayLine      : string := "";		-- "0_to_63_delay_value"
    outputCapacity       : string := "";		-- 0 to 40 (value in pF)
    -- Delay Control
    spath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay

);
port (
    FCK	: in std_logic := '0';
    SCK	: in std_logic := '0';
    R	: in std_logic := '0';
    I	: in std_logic_vector(data_size - 1 downto 0) := (others => '0');
    IO	: out std_logic := '0';
    -- Delay Control
    DCK	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DS	: in std_logic_vector(1 downto 0) := (others => '0');
    DRA	: in std_logic_vector(5 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');
    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0')
);
end component NX_SER;

component NX_DES is
generic (
    data_size            : integer range 2 to 10 := 5;	-- -- Pad location Number of deserialization factor
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0") or differential ("1")
    termination          : string := "";		-- Input impedance adaptatio    terminationReference : string := "";
    terminationReference : string := "";		-- "floating" or "VTT"
    turbo                : string := "";		-- Input impedance adaptation
    weakTermination      : string := "";		-- "floating" or "VTT"
    inputDelayLine       : string := "";		-- "0_to_63_delay_value"
    inputSignalSlope     : string := "";		-- Decimal value "0.5" to "20" (value in V/ns)
    -- Delay Control
    dpath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay

);
port (
    FCK	: in std_logic := '0';
    SCK	: in std_logic := '0';
    R	: in std_logic := '0';
    IO	: in std_logic := '0';
    O	: out std_logic_vector(data_size - 1 downto 0) := (others => '0');
    -- Delay Control
    DCK	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DS	: in std_logic_vector(1 downto 0) := (others => '0');
    DRA	: in std_logic_vector(5 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');
    FZ	: in std_logic := '0';
    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0');
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0'
);
end component NX_DES;

component NX_SERDES is
generic (
    data_size            : integer range 2 to 10 := 5;	-- Serialiser/deserializer factor 
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0" or differential ("1")
    slewRate             : string := "";		-- Slow, Medium or Fast
    termination          : string := "";		-- Input impedance adaptation
    terminationReference : string := "";		-- "floating" or "VTT"
    turbo                : string := "";		-- "true" or "false"
    weakTermination      : string := "";		-- "PullUp" or "None"
    inputDelayLine       : string := "";		-- "O_to_63_delay_value"
    outputDelayLine      : string := "";		-- "O_to_63_delay_value"
    inputSignalSlope     : string := "";		-- Decimal value "0.5" to "20" (value in V/ns)
    outputCapacity       : string := "";		-- "0" to "40" (value in pF)
    cpath_registered     : bit := '0';			-- Use Register in Enable Path ('1')
    -- Delay Control
    spath_dynamic        : bit := '0';			-- 0: off/fixed delay, 1: dynamic delay
    dpath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay
);
port (
    FCK	: in std_logic := '0';
    SCK	: in std_logic := '0';
    RTX	: in std_logic := '0';
    RRX	: in std_logic := '0';
    CI	: in std_logic := '0';
    CCK	: in std_logic := '0';
    CL	: in std_logic := '0';
    CR	: in std_logic := '0';
    I	: in std_logic_vector(data_size - 1 downto 0) := (others => '0');
    IO	: inout std_logic := '0';
    O	: out std_logic_vector(data_size - 1 downto 0) := (others => '0');
    -- Delay Control
    DCK	: in std_logic := '0';
    DRL	: in std_logic := '0';
    DIG	: in std_logic := '0';
    DS	: in std_logic_vector(1 downto 0) := (others => '0');
    DRA	: in std_logic_vector(5 downto 0) := (others => '0');
    DRI	: in std_logic_vector(5 downto 0) := (others => '0');
    FZ	: in std_logic := '0';
    DRO	: out std_logic_vector(5 downto 0) := (others => '0');
    DID	: out std_logic_vector(5 downto 0) := (others => '0');
    FLD	: out std_logic := '0';
    FLG	: out std_logic := '0'
);
end component NX_SERDES;

component NX_SERVICE_U is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    fabric_otp_user_tst_scanenable_i	: in std_logic := '0';
    fabric_otp_cfg_loader_read_en_i	: in std_logic := '0';
    fabric_otp_security_force_pdn1_i	: in std_logic := '0';
    fabric_otp_security_scanenable_i	: in std_logic := '0';
    fabric_otp_user_din_i1	: in std_logic := '0';
    fabric_otp_user_din_i2	: in std_logic := '0';
    fabric_otp_user_din_i3	: in std_logic := '0';
    fabric_otp_user_din_i4	: in std_logic := '0';
    fabric_otp_user_din_i5	: in std_logic := '0';
    fabric_otp_user_din_i6	: in std_logic := '0';
    fabric_otp_user_din_i7	: in std_logic := '0';
    fabric_otp_user_din_i8	: in std_logic := '0';
    fabric_otp_user_din_i9	: in std_logic := '0';
    fabric_otp_user_din_i10	: in std_logic := '0';
    fabric_otp_user_din_i11	: in std_logic := '0';
    fabric_otp_user_din_i12	: in std_logic := '0';
    fabric_otp_user_din_i13	: in std_logic := '0';
    fabric_otp_user_din_i14	: in std_logic := '0';
    fabric_otp_user_din_i15	: in std_logic := '0';
    fabric_otp_user_din_i16	: in std_logic := '0';
    fabric_otp_user_din_i17	: in std_logic := '0';
    fabric_otp_user_din_i18	: in std_logic := '0';
    fabric_otp_user_din_i19	: in std_logic := '0';
    fabric_otp_user_din_i20	: in std_logic := '0';
    fabric_otp_user_din_i21	: in std_logic := '0';
    fabric_otp_user_din_i22	: in std_logic := '0';
    fabric_otp_user_din_i23	: in std_logic := '0';
    fabric_otp_user_din_i24	: in std_logic := '0';
    fabric_otp_user_din_i25	: in std_logic := '0';
    fabric_otp_user_din_i26	: in std_logic := '0';
    fabric_otp_user_din_i27	: in std_logic := '0';
    fabric_otp_user_din_i28	: in std_logic := '0';
    fabric_otp_user_din_i29	: in std_logic := '0';
    fabric_otp_user_din_i30	: in std_logic := '0';
    fabric_otp_user_din_i31	: in std_logic := '0';
    fabric_otp_user_din_i32	: in std_logic := '0';
    fabric_otp_user_din_i33	: in std_logic := '0';
    fabric_otp_user_din_i34	: in std_logic := '0';
    fabric_otp_user_din_i35	: in std_logic := '0';
    fabric_otp_user_din_i36	: in std_logic := '0';
    fabric_otp_user_din_i37	: in std_logic := '0';
    fabric_otp_user_din_i38	: in std_logic := '0';
    fabric_otp_user_din_i39	: in std_logic := '0';
    fabric_mrepair_fuse_prgwidth_i1	: in std_logic := '0';
    fabric_mrepair_fuse_prgwidth_i2	: in std_logic := '0';
    fabric_mrepair_fuse_prgwidth_i3	: in std_logic := '0';
    fabric_otp_apb_wdata_i1	: in std_logic := '0';
    fabric_otp_apb_wdata_i2	: in std_logic := '0';
    fabric_otp_apb_wdata_i3	: in std_logic := '0';
    fabric_otp_apb_wdata_i4	: in std_logic := '0';
    fabric_otp_apb_wdata_i5	: in std_logic := '0';
    fabric_otp_apb_wdata_i6	: in std_logic := '0';
    fabric_otp_apb_wdata_i7	: in std_logic := '0';
    fabric_otp_apb_wdata_i8	: in std_logic := '0';
    fabric_otp_apb_wdata_i9	: in std_logic := '0';
    fabric_otp_apb_wdata_i10	: in std_logic := '0';
    fabric_otp_apb_wdata_i11	: in std_logic := '0';
    fabric_otp_apb_wdata_i12	: in std_logic := '0';
    fabric_otp_apb_wdata_i13	: in std_logic := '0';
    fabric_otp_apb_wdata_i14	: in std_logic := '0';
    fabric_otp_apb_wdata_i15	: in std_logic := '0';
    fabric_otp_apb_wdata_i16	: in std_logic := '0';
    fabric_otp_apb_wdata_i17	: in std_logic := '0';
    fabric_otp_apb_wdata_i18	: in std_logic := '0';
    fabric_otp_apb_wdata_i19	: in std_logic := '0';
    fabric_otp_apb_wdata_i20	: in std_logic := '0';
    fabric_otp_apb_wdata_i21	: in std_logic := '0';
    fabric_otp_apb_wdata_i22	: in std_logic := '0';
    fabric_otp_apb_wdata_i23	: in std_logic := '0';
    fabric_otp_apb_wdata_i24	: in std_logic := '0';
    fabric_otp_apb_wdata_i25	: in std_logic := '0';
    fabric_otp_apb_wdata_i26	: in std_logic := '0';
    fabric_otp_apb_wdata_i27	: in std_logic := '0';
    fabric_otp_apb_wdata_i28	: in std_logic := '0';
    fabric_otp_apb_wdata_i29	: in std_logic := '0';
    fabric_otp_apb_wdata_i30	: in std_logic := '0';
    fabric_otp_apb_wdata_i31	: in std_logic := '0';
    fabric_otp_apb_wdata_i32	: in std_logic := '0';
    fabric_otp_cfg_clk_otpm_disable_i	: in std_logic := '0';
    fabric_otp_user_disturbcheck_i	: in std_logic := '0';
    fabric_mrepair_fuse_read_i	: in std_logic := '0';
    fabric_otp_user_rbact2_i	: in std_logic := '0';
    fabric_mrepair_fuse_eccbypass_i	: in std_logic := '0';
    fabric_otp_user_bistmode_i	: in std_logic := '0';
    fabric_otp_user_add_i1	: in std_logic := '0';
    fabric_otp_user_add_i2	: in std_logic := '0';
    fabric_otp_user_add_i3	: in std_logic := '0';
    fabric_otp_user_add_i4	: in std_logic := '0';
    fabric_otp_user_add_i5	: in std_logic := '0';
    fabric_otp_user_add_i6	: in std_logic := '0';
    fabric_otp_user_add_i7	: in std_logic := '0';
    fabric_otp_user_tm_i	: in std_logic := '0';
    fabric_otp_rstn_i	: in std_logic := '0';
    fabric_mrepair_fuse_disturbchecked_i	: in std_logic := '0';
    fabric_otp_user_rbact1_i	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i1	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i2	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i3	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i4	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i5	: in std_logic := '0';
    fabric_parusr_type_i1	: in std_logic := '0';
    fabric_parusr_type_i2	: in std_logic := '0';
    fabric_mrepair_fuse_redbypass_i	: in std_logic := '0';
    fabric_otp_user_eccbypass_i	: in std_logic := '0';
    fabric_otp_user_redbypass_i	: in std_logic := '0';
    fabric_mrepair_mode_i1	: in std_logic := '0';
    fabric_mrepair_mode_i2	: in std_logic := '0';
    fabric_mrepair_mode_i3	: in std_logic := '0';
    fabric_mrepair_mode_i4	: in std_logic := '0';
    fabric_parusr_cs_i	: in std_logic := '0';
    fabric_sif_reg_en_i1	: in std_logic := '0';
    fabric_sif_reg_en_i2	: in std_logic := '0';
    fabric_sif_reg_en_i3	: in std_logic := '0';
    fabric_sif_reg_en_i4	: in std_logic := '0';
    fabric_sif_reg_en_i5	: in std_logic := '0';
    fabric_sif_reg_en_i6	: in std_logic := '0';
    fabric_sif_reg_en_i7	: in std_logic := '0';
    fabric_sif_reg_en_i8	: in std_logic := '0';
    fabric_sif_reg_en_i9	: in std_logic := '0';
    fabric_sif_reg_en_i10	: in std_logic := '0';
    fabric_sif_reg_en_i11	: in std_logic := '0';
    fabric_sif_reg_en_i12	: in std_logic := '0';
    fabric_sif_reg_en_i13	: in std_logic := '0';
    fabric_sif_reg_en_i14	: in std_logic := '0';
    fabric_sif_reg_en_i15	: in std_logic := '0';
    fabric_sif_reg_en_i16	: in std_logic := '0';
    fabric_sif_reg_en_i17	: in std_logic := '0';
    fabric_sif_reg_en_i18	: in std_logic := '0';
    fabric_sif_reg_en_i19	: in std_logic := '0';
    fabric_sif_reg_en_i20	: in std_logic := '0';
    fabric_sif_reg_en_i21	: in std_logic := '0';
    fabric_sif_reg_en_i22	: in std_logic := '0';
    fabric_sif_reg_en_i23	: in std_logic := '0';
    fabric_sif_reg_en_i24	: in std_logic := '0';
    fabric_sif_reg_en_i25	: in std_logic := '0';
    fabric_sif_reg_en_i26	: in std_logic := '0';
    fabric_sif_reg_en_i27	: in std_logic := '0';
    fabric_sif_reg_en_i28	: in std_logic := '0';
    fabric_sif_reg_en_i29	: in std_logic := '0';
    fabric_sif_reg_en_i30	: in std_logic := '0';
    fabric_sif_reg_en_i31	: in std_logic := '0';
    fabric_sif_reg_en_i32	: in std_logic := '0';
    fabric_sif_reg_en_i33	: in std_logic := '0';
    fabric_sif_reg_en_i34	: in std_logic := '0';
    fabric_sif_reg_en_i35	: in std_logic := '0';
    fabric_sif_reg_en_i36	: in std_logic := '0';
    fabric_sif_reg_en_i37	: in std_logic := '0';
    fabric_sif_reg_en_i38	: in std_logic := '0';
    fabric_sif_reg_en_i39	: in std_logic := '0';
    fabric_sif_reg_en_i40	: in std_logic := '0';
    fabric_sif_reg_en_i41	: in std_logic := '0';
    fabric_sif_reg_en_i42	: in std_logic := '0';
    fabric_sif_reg_en_i43	: in std_logic := '0';
    fabric_sif_reg_en_i44	: in std_logic := '0';
    fabric_sif_reg_en_i45	: in std_logic := '0';
    fabric_sif_reg_en_i46	: in std_logic := '0';
    fabric_sif_reg_en_i47	: in std_logic := '0';
    fabric_sif_reg_en_i48	: in std_logic := '0';
    fabric_sif_reg_en_i49	: in std_logic := '0';
    fabric_sif_reg_en_i50	: in std_logic := '0';
    fabric_sif_reg_en_i51	: in std_logic := '0';
    fabric_sif_reg_en_i52	: in std_logic := '0';
    fabric_sif_reg_en_i53	: in std_logic := '0';
    fabric_sif_reg_en_i54	: in std_logic := '0';
    fabric_sif_reg_en_i55	: in std_logic := '0';
    fabric_sif_reg_en_i56	: in std_logic := '0';
    fabric_sif_reg_en_i57	: in std_logic := '0';
    fabric_sif_reg_en_i58	: in std_logic := '0';
    fabric_sif_reg_en_i59	: in std_logic := '0';
    fabric_sif_reg_en_i60	: in std_logic := '0';
    fabric_sif_reg_en_i61	: in std_logic := '0';
    fabric_sif_reg_en_i62	: in std_logic := '0';
    fabric_sif_reg_en_i63	: in std_logic := '0';
    fabric_sif_reg_en_i64	: in std_logic := '0';
    fabric_sif_reg_en_i65	: in std_logic := '0';
    fabric_sif_reg_en_i66	: in std_logic := '0';
    fabric_sif_reg_en_i67	: in std_logic := '0';
    fabric_sif_reg_en_i68	: in std_logic := '0';
    fabric_sif_reg_en_i69	: in std_logic := '0';
    fabric_sif_reg_en_i70	: in std_logic := '0';
    fabric_sif_reg_en_i71	: in std_logic := '0';
    fabric_sif_reg_en_i72	: in std_logic := '0';
    fabric_sif_reg_en_i73	: in std_logic := '0';
    fabric_sif_reg_en_i74	: in std_logic := '0';
    fabric_sif_reg_en_i75	: in std_logic := '0';
    fabric_sif_reg_en_i76	: in std_logic := '0';
    fabric_sif_reg_en_i77	: in std_logic := '0';
    fabric_sif_reg_en_i78	: in std_logic := '0';
    fabric_sif_reg_en_i79	: in std_logic := '0';
    fabric_sif_reg_en_i80	: in std_logic := '0';
    fabric_sif_reg_en_i81	: in std_logic := '0';
    fabric_sif_reg_en_i82	: in std_logic := '0';
    fabric_sif_reg_en_i83	: in std_logic := '0';
    fabric_sif_reg_en_i84	: in std_logic := '0';
    fabric_sif_reg_en_i85	: in std_logic := '0';
    fabric_sif_reg_en_i86	: in std_logic := '0';
    fabric_sif_reg_en_i87	: in std_logic := '0';
    fabric_sif_reg_en_i88	: in std_logic := '0';
    fabric_sif_reg_en_i89	: in std_logic := '0';
    fabric_sif_reg_en_i90	: in std_logic := '0';
    fabric_sif_reg_en_i91	: in std_logic := '0';
    fabric_sif_reg_en_i92	: in std_logic := '0';
    fabric_sif_reg_en_i93	: in std_logic := '0';
    fabric_sif_reg_en_i94	: in std_logic := '0';
    fabric_sif_reg_en_i95	: in std_logic := '0';
    fabric_sif_reg_en_i96	: in std_logic := '0';
    fabric_sif_reg_en_i97	: in std_logic := '0';
    fabric_sif_reg_en_i98	: in std_logic := '0';
    fabric_sif_reg_en_i99	: in std_logic := '0';
    fabric_sif_reg_en_i100	: in std_logic := '0';
    fabric_sif_reg_en_i101	: in std_logic := '0';
    fabric_sif_reg_en_i102	: in std_logic := '0';
    fabric_sif_reg_en_i103	: in std_logic := '0';
    fabric_sif_reg_en_i104	: in std_logic := '0';
    fabric_sif_reg_en_i105	: in std_logic := '0';
    fabric_sif_reg_en_i106	: in std_logic := '0';
    fabric_sif_reg_en_i107	: in std_logic := '0';
    fabric_sif_reg_en_i108	: in std_logic := '0';
    fabric_sif_reg_en_i109	: in std_logic := '0';
    fabric_sif_reg_en_i110	: in std_logic := '0';
    fabric_sif_reg_en_i111	: in std_logic := '0';
    fabric_sif_reg_en_i112	: in std_logic := '0';
    fabric_sif_reg_en_i113	: in std_logic := '0';
    fabric_sif_reg_en_i114	: in std_logic := '0';
    fabric_sif_reg_en_i115	: in std_logic := '0';
    fabric_sif_reg_en_i116	: in std_logic := '0';
    fabric_sif_reg_en_i117	: in std_logic := '0';
    fabric_sif_reg_en_i118	: in std_logic := '0';
    fabric_sif_reg_en_i119	: in std_logic := '0';
    fabric_sif_reg_en_i120	: in std_logic := '0';
    fabric_mrepair_fuse_rbact2_i	: in std_logic := '0';
    fabric_data_from_system_i	: in std_logic := '0';
    fabric_data_from_bist_i1	: in std_logic := '0';
    fabric_data_from_bist_i2	: in std_logic := '0';
    fabric_data_from_bist_i3	: in std_logic := '0';
    fabric_data_from_bist_i4	: in std_logic := '0';
    fabric_data_from_bist_i5	: in std_logic := '0';
    fabric_data_from_bist_i6	: in std_logic := '0';
    fabric_data_from_bist_i7	: in std_logic := '0';
    fabric_data_from_bist_i8	: in std_logic := '0';
    fabric_data_from_bist_i9	: in std_logic := '0';
    fabric_data_from_bist_i10	: in std_logic := '0';
    fabric_data_from_bist_i11	: in std_logic := '0';
    fabric_data_from_bist_i12	: in std_logic := '0';
    fabric_data_from_bist_i13	: in std_logic := '0';
    fabric_data_from_bist_i14	: in std_logic := '0';
    fabric_data_from_bist_i15	: in std_logic := '0';
    fabric_data_from_bist_i16	: in std_logic := '0';
    fabric_data_from_bist_i17	: in std_logic := '0';
    fabric_data_from_bist_i18	: in std_logic := '0';
    fabric_data_from_bist_i19	: in std_logic := '0';
    fabric_data_from_bist_i20	: in std_logic := '0';
    fabric_data_from_bist_i21	: in std_logic := '0';
    fabric_data_from_bist_i22	: in std_logic := '0';
    fabric_data_from_bist_i23	: in std_logic := '0';
    fabric_data_from_bist_i24	: in std_logic := '0';
    fabric_otp_apb_enable_i	: in std_logic := '0';
    fabric_mrepair_fuse_tm_i	: in std_logic := '0';
    fabric_otp_security_rbact2_i	: in std_logic := '0';
    fabric_otp_security_rbact1_i	: in std_logic := '0';
    fabric_shift_en_i1	: in std_logic := '0';
    fabric_shift_en_i2	: in std_logic := '0';
    fabric_shift_en_i3	: in std_logic := '0';
    fabric_shift_en_i4	: in std_logic := '0';
    fabric_shift_en_i5	: in std_logic := '0';
    fabric_shift_en_i6	: in std_logic := '0';
    fabric_shift_en_i7	: in std_logic := '0';
    fabric_shift_en_i8	: in std_logic := '0';
    fabric_shift_en_i9	: in std_logic := '0';
    fabric_shift_en_i10	: in std_logic := '0';
    fabric_shift_en_i11	: in std_logic := '0';
    fabric_shift_en_i12	: in std_logic := '0';
    fabric_shift_en_i13	: in std_logic := '0';
    fabric_shift_en_i14	: in std_logic := '0';
    fabric_shift_en_i15	: in std_logic := '0';
    fabric_shift_en_i16	: in std_logic := '0';
    fabric_shift_en_i17	: in std_logic := '0';
    fabric_shift_en_i18	: in std_logic := '0';
    fabric_shift_en_i19	: in std_logic := '0';
    fabric_shift_en_i20	: in std_logic := '0';
    fabric_shift_en_i21	: in std_logic := '0';
    fabric_shift_en_i22	: in std_logic := '0';
    fabric_shift_en_i23	: in std_logic := '0';
    fabric_shift_en_i24	: in std_logic := '0';
    fabric_otp_cfg_loader_write_en_i	: in std_logic := '0';
    fabric_user_data_i1	: in std_logic := '0';
    fabric_user_data_i2	: in std_logic := '0';
    fabric_user_data_i3	: in std_logic := '0';
    fabric_user_data_i4	: in std_logic := '0';
    fabric_user_data_i5	: in std_logic := '0';
    fabric_user_data_i6	: in std_logic := '0';
    fabric_user_data_i7	: in std_logic := '0';
    fabric_user_data_i8	: in std_logic := '0';
    fabric_user_data_i9	: in std_logic := '0';
    fabric_user_data_i10	: in std_logic := '0';
    fabric_user_data_i11	: in std_logic := '0';
    fabric_user_data_i12	: in std_logic := '0';
    fabric_user_data_i13	: in std_logic := '0';
    fabric_user_data_i14	: in std_logic := '0';
    fabric_user_data_i15	: in std_logic := '0';
    fabric_user_data_i16	: in std_logic := '0';
    fabric_user_data_i17	: in std_logic := '0';
    fabric_user_data_i18	: in std_logic := '0';
    fabric_user_data_i19	: in std_logic := '0';
    fabric_user_data_i20	: in std_logic := '0';
    fabric_user_data_i21	: in std_logic := '0';
    fabric_user_data_i22	: in std_logic := '0';
    fabric_user_data_i23	: in std_logic := '0';
    fabric_user_data_i24	: in std_logic := '0';
    fabric_user_data_i25	: in std_logic := '0';
    fabric_user_data_i26	: in std_logic := '0';
    fabric_user_data_i27	: in std_logic := '0';
    fabric_user_data_i28	: in std_logic := '0';
    fabric_user_data_i29	: in std_logic := '0';
    fabric_user_data_i30	: in std_logic := '0';
    fabric_user_data_i31	: in std_logic := '0';
    fabric_user_data_i32	: in std_logic := '0';
    fabric_mrepair_fuse_suppadd_i	: in std_logic := '0';
    fabric_mrepair_fuse_prog_i	: in std_logic := '0';
    fabric_otp_user_wordlock_i	: in std_logic := '0';
    fabric_ahb_direct_data_i1	: in std_logic := '0';
    fabric_ahb_direct_data_i2	: in std_logic := '0';
    fabric_ahb_direct_data_i3	: in std_logic := '0';
    fabric_ahb_direct_data_i4	: in std_logic := '0';
    fabric_ahb_direct_data_i5	: in std_logic := '0';
    fabric_ahb_direct_data_i6	: in std_logic := '0';
    fabric_ahb_direct_data_i7	: in std_logic := '0';
    fabric_ahb_direct_data_i8	: in std_logic := '0';
    fabric_ahb_direct_data_i9	: in std_logic := '0';
    fabric_ahb_direct_data_i10	: in std_logic := '0';
    fabric_ahb_direct_data_i11	: in std_logic := '0';
    fabric_ahb_direct_data_i12	: in std_logic := '0';
    fabric_ahb_direct_data_i13	: in std_logic := '0';
    fabric_ahb_direct_data_i14	: in std_logic := '0';
    fabric_ahb_direct_data_i15	: in std_logic := '0';
    fabric_ahb_direct_data_i16	: in std_logic := '0';
    fabric_ahb_direct_data_i17	: in std_logic := '0';
    fabric_ahb_direct_data_i18	: in std_logic := '0';
    fabric_ahb_direct_data_i19	: in std_logic := '0';
    fabric_ahb_direct_data_i20	: in std_logic := '0';
    fabric_ahb_direct_data_i21	: in std_logic := '0';
    fabric_ahb_direct_data_i22	: in std_logic := '0';
    fabric_ahb_direct_data_i23	: in std_logic := '0';
    fabric_ahb_direct_data_i24	: in std_logic := '0';
    fabric_ahb_direct_data_i25	: in std_logic := '0';
    fabric_ahb_direct_data_i26	: in std_logic := '0';
    fabric_ahb_direct_data_i27	: in std_logic := '0';
    fabric_ahb_direct_data_i28	: in std_logic := '0';
    fabric_ahb_direct_data_i29	: in std_logic := '0';
    fabric_ahb_direct_data_i30	: in std_logic := '0';
    fabric_ahb_direct_data_i31	: in std_logic := '0';
    fabric_ahb_direct_data_i32	: in std_logic := '0';
    fabric_otp_user_prog_i	: in std_logic := '0';
    fabric_pd_active_i1	: in std_logic := '0';
    fabric_pd_active_i2	: in std_logic := '0';
    fabric_pd_active_i3	: in std_logic := '0';
    fabric_pd_active_i4	: in std_logic := '0';
    fabric_pd_active_i5	: in std_logic := '0';
    fabric_pd_active_i6	: in std_logic := '0';
    fabric_pd_active_i7	: in std_logic := '0';
    fabric_pd_active_i8	: in std_logic := '0';
    fabric_pd_active_i9	: in std_logic := '0';
    fabric_pd_active_i10	: in std_logic := '0';
    fabric_pd_active_i11	: in std_logic := '0';
    fabric_pd_active_i12	: in std_logic := '0';
    fabric_pd_active_i13	: in std_logic := '0';
    fabric_pd_active_i14	: in std_logic := '0';
    fabric_pd_active_i15	: in std_logic := '0';
    fabric_pd_active_i16	: in std_logic := '0';
    fabric_pd_active_i17	: in std_logic := '0';
    fabric_pd_active_i18	: in std_logic := '0';
    fabric_pd_active_i19	: in std_logic := '0';
    fabric_pd_active_i20	: in std_logic := '0';
    fabric_pd_active_i21	: in std_logic := '0';
    fabric_pd_active_i22	: in std_logic := '0';
    fabric_pd_active_i23	: in std_logic := '0';
    fabric_pd_active_i24	: in std_logic := '0';
    fabric_otp_user_suppadd_i	: in std_logic := '0';
    fabric_mrepair_fuse_pdn_i	: in std_logic := '0';
    fabric_otp_security_scanin_i1	: in std_logic := '0';
    fabric_otp_security_scanin_i2	: in std_logic := '0';
    fabric_otp_security_scanin_i3	: in std_logic := '0';
    fabric_otp_security_scanin_i4	: in std_logic := '0';
    fabric_otp_security_scanin_i5	: in std_logic := '0';
    fabric_end_encoding_i	: in std_logic := '0';
    fabric_jtag_tdo_usr2_i	: in std_logic := '0';
    fabric_mrepair_fuse_wordlock_i	: in std_logic := '0';
    fabric_otp_user_prgwidth_i1	: in std_logic := '0';
    fabric_otp_user_prgwidth_i2	: in std_logic := '0';
    fabric_otp_user_prgwidth_i3	: in std_logic := '0';
    fabric_otp_user_read_i	: in std_logic := '0';
    fabric_mrepair_fuse_add_i1	: in std_logic := '0';
    fabric_mrepair_fuse_add_i2	: in std_logic := '0';
    fabric_mrepair_fuse_add_i3	: in std_logic := '0';
    fabric_mrepair_fuse_add_i4	: in std_logic := '0';
    fabric_mrepair_fuse_add_i5	: in std_logic := '0';
    fabric_mrepair_fuse_add_i6	: in std_logic := '0';
    fabric_mrepair_fuse_add_i7	: in std_logic := '0';
    fabric_mrepair_fuse_bistmode_i	: in std_logic := '0';
    fabric_jtag_tdo_usr1_i	: in std_logic := '0';
    fabric_otp_cfg_clk_fab_en_i	: in std_logic := '0';
    fabric_io_in_i1	: in std_logic := '0';
    fabric_io_in_i2	: in std_logic := '0';
    fabric_io_in_i3	: in std_logic := '0';
    fabric_io_in_i4	: in std_logic := '0';
    fabric_io_in_i5	: in std_logic := '0';
    fabric_io_in_i6	: in std_logic := '0';
    fabric_io_in_i7	: in std_logic := '0';
    fabric_io_in_i8	: in std_logic := '0';
    fabric_io_in_i9	: in std_logic := '0';
    fabric_io_in_i10	: in std_logic := '0';
    fabric_io_in_i11	: in std_logic := '0';
    fabric_io_in_i12	: in std_logic := '0';
    fabric_io_in_i13	: in std_logic := '0';
    fabric_io_in_i14	: in std_logic := '0';
    fabric_io_in_i15	: in std_logic := '0';
    fabric_io_in_i16	: in std_logic := '0';
    fabric_io_in_i17	: in std_logic := '0';
    fabric_io_in_i18	: in std_logic := '0';
    fabric_io_in_i19	: in std_logic := '0';
    fabric_io_in_i20	: in std_logic := '0';
    fabric_io_in_i21	: in std_logic := '0';
    fabric_io_in_i22	: in std_logic := '0';
    fabric_io_in_i23	: in std_logic := '0';
    fabric_io_in_i24	: in std_logic := '0';
    fabric_io_in_i25	: in std_logic := '0';
    fabric_sif_load_en_i1	: in std_logic := '0';
    fabric_sif_load_en_i2	: in std_logic := '0';
    fabric_sif_load_en_i3	: in std_logic := '0';
    fabric_sif_load_en_i4	: in std_logic := '0';
    fabric_sif_load_en_i5	: in std_logic := '0';
    fabric_sif_load_en_i6	: in std_logic := '0';
    fabric_sif_load_en_i7	: in std_logic := '0';
    fabric_sif_load_en_i8	: in std_logic := '0';
    fabric_sif_load_en_i9	: in std_logic := '0';
    fabric_sif_load_en_i10	: in std_logic := '0';
    fabric_sif_load_en_i11	: in std_logic := '0';
    fabric_sif_load_en_i12	: in std_logic := '0';
    fabric_sif_load_en_i13	: in std_logic := '0';
    fabric_sif_load_en_i14	: in std_logic := '0';
    fabric_sif_load_en_i15	: in std_logic := '0';
    fabric_sif_load_en_i16	: in std_logic := '0';
    fabric_sif_load_en_i17	: in std_logic := '0';
    fabric_sif_load_en_i18	: in std_logic := '0';
    fabric_sif_load_en_i19	: in std_logic := '0';
    fabric_sif_load_en_i20	: in std_logic := '0';
    fabric_sif_load_en_i21	: in std_logic := '0';
    fabric_sif_load_en_i22	: in std_logic := '0';
    fabric_sif_load_en_i23	: in std_logic := '0';
    fabric_sif_load_en_i24	: in std_logic := '0';
    fabric_mrepair_fuse_din_i1	: in std_logic := '0';
    fabric_mrepair_fuse_din_i2	: in std_logic := '0';
    fabric_mrepair_fuse_din_i3	: in std_logic := '0';
    fabric_mrepair_fuse_din_i4	: in std_logic := '0';
    fabric_mrepair_fuse_din_i5	: in std_logic := '0';
    fabric_mrepair_fuse_din_i6	: in std_logic := '0';
    fabric_mrepair_fuse_din_i7	: in std_logic := '0';
    fabric_mrepair_fuse_din_i8	: in std_logic := '0';
    fabric_mrepair_fuse_din_i9	: in std_logic := '0';
    fabric_mrepair_fuse_din_i10	: in std_logic := '0';
    fabric_mrepair_fuse_din_i11	: in std_logic := '0';
    fabric_mrepair_fuse_din_i12	: in std_logic := '0';
    fabric_mrepair_fuse_din_i13	: in std_logic := '0';
    fabric_mrepair_fuse_din_i14	: in std_logic := '0';
    fabric_mrepair_fuse_din_i15	: in std_logic := '0';
    fabric_mrepair_fuse_din_i16	: in std_logic := '0';
    fabric_mrepair_fuse_din_i17	: in std_logic := '0';
    fabric_mrepair_fuse_din_i18	: in std_logic := '0';
    fabric_mrepair_fuse_din_i19	: in std_logic := '0';
    fabric_mrepair_fuse_din_i20	: in std_logic := '0';
    fabric_mrepair_fuse_din_i21	: in std_logic := '0';
    fabric_mrepair_fuse_din_i22	: in std_logic := '0';
    fabric_mrepair_fuse_din_i23	: in std_logic := '0';
    fabric_mrepair_fuse_din_i24	: in std_logic := '0';
    fabric_mrepair_fuse_din_i25	: in std_logic := '0';
    fabric_mrepair_fuse_din_i26	: in std_logic := '0';
    fabric_mrepair_fuse_din_i27	: in std_logic := '0';
    fabric_mrepair_fuse_din_i28	: in std_logic := '0';
    fabric_mrepair_fuse_din_i29	: in std_logic := '0';
    fabric_mrepair_fuse_din_i30	: in std_logic := '0';
    fabric_mrepair_fuse_din_i31	: in std_logic := '0';
    fabric_mrepair_fuse_din_i32	: in std_logic := '0';
    fabric_mrepair_fuse_din_i33	: in std_logic := '0';
    fabric_mrepair_fuse_din_i34	: in std_logic := '0';
    fabric_mrepair_fuse_din_i35	: in std_logic := '0';
    fabric_mrepair_fuse_din_i36	: in std_logic := '0';
    fabric_mrepair_fuse_din_i37	: in std_logic := '0';
    fabric_mrepair_fuse_din_i38	: in std_logic := '0';
    fabric_mrepair_fuse_din_i39	: in std_logic := '0';
    fabric_otp_apb_addr_i1	: in std_logic := '0';
    fabric_otp_apb_addr_i2	: in std_logic := '0';
    fabric_otp_apb_addr_i3	: in std_logic := '0';
    fabric_otp_apb_addr_i4	: in std_logic := '0';
    fabric_otp_apb_addr_i5	: in std_logic := '0';
    fabric_otp_apb_addr_i6	: in std_logic := '0';
    fabric_otp_apb_addr_i7	: in std_logic := '0';
    fabric_otp_apb_addr_i8	: in std_logic := '0';
    fabric_otp_apb_addr_i9	: in std_logic := '0';
    fabric_otp_apb_addr_i10	: in std_logic := '0';
    fabric_otp_apb_addr_i11	: in std_logic := '0';
    fabric_otp_apb_addr_i12	: in std_logic := '0';
    fabric_otp_apb_addr_i13	: in std_logic := '0';
    fabric_otp_apb_addr_i14	: in std_logic := '0';
    fabric_otp_apb_addr_i15	: in std_logic := '0';
    fabric_otp_apb_addr_i16	: in std_logic := '0';
    fabric_otp_apb_addr_i17	: in std_logic := '0';
    fabric_otp_apb_addr_i18	: in std_logic := '0';
    fabric_otp_apb_addr_i19	: in std_logic := '0';
    fabric_otp_apb_addr_i20	: in std_logic := '0';
    fabric_otp_apb_addr_i21	: in std_logic := '0';
    fabric_otp_apb_addr_i22	: in std_logic := '0';
    fabric_otp_apb_addr_i23	: in std_logic := '0';
    fabric_otp_apb_addr_i24	: in std_logic := '0';
    fabric_otp_apb_addr_i25	: in std_logic := '0';
    fabric_otp_apb_addr_i26	: in std_logic := '0';
    fabric_otp_apb_addr_i27	: in std_logic := '0';
    fabric_otp_apb_addr_i28	: in std_logic := '0';
    fabric_otp_apb_addr_i29	: in std_logic := '0';
    fabric_otp_apb_addr_i30	: in std_logic := '0';
    fabric_otp_apb_addr_i31	: in std_logic := '0';
    fabric_otp_apb_addr_i32	: in std_logic := '0';
    fabric_otp_apb_sel_i	: in std_logic := '0';
    fabric_mrepair_fuse_rbact1_i	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i1	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i2	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i3	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i4	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i5	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i6	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i7	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i8	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i9	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i10	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i11	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i12	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i13	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i14	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i15	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i16	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i17	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i18	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i19	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i20	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i21	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i22	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i23	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i24	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i25	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i26	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i27	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i28	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i29	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i30	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i31	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i32	: in std_logic := '0';
    fabric_otp_cfg_fabric_apb_en_i	: in std_logic := '0';
    fabric_data_shift_en_i	: in std_logic := '0';
    fabric_lowskew_i21	: in std_logic := '0';
    fabric_direct_data_i1	: in std_logic := '0';
    fabric_direct_data_i2	: in std_logic := '0';
    fabric_direct_data_i3	: in std_logic := '0';
    fabric_direct_data_i4	: in std_logic := '0';
    fabric_direct_data_i5	: in std_logic := '0';
    fabric_direct_data_i6	: in std_logic := '0';
    fabric_direct_data_i7	: in std_logic := '0';
    fabric_direct_data_i8	: in std_logic := '0';
    fabric_direct_data_i9	: in std_logic := '0';
    fabric_direct_data_i10	: in std_logic := '0';
    fabric_direct_data_i11	: in std_logic := '0';
    fabric_direct_data_i12	: in std_logic := '0';
    fabric_direct_data_i13	: in std_logic := '0';
    fabric_direct_data_i14	: in std_logic := '0';
    fabric_direct_data_i15	: in std_logic := '0';
    fabric_direct_data_i16	: in std_logic := '0';
    fabric_direct_data_i17	: in std_logic := '0';
    fabric_direct_data_i18	: in std_logic := '0';
    fabric_direct_data_i19	: in std_logic := '0';
    fabric_direct_data_i20	: in std_logic := '0';
    fabric_direct_data_i21	: in std_logic := '0';
    fabric_direct_data_i22	: in std_logic := '0';
    fabric_direct_data_i23	: in std_logic := '0';
    fabric_direct_data_i24	: in std_logic := '0';
    fabric_direct_data_i25	: in std_logic := '0';
    fabric_direct_data_i26	: in std_logic := '0';
    fabric_direct_data_i27	: in std_logic := '0';
    fabric_direct_data_i28	: in std_logic := '0';
    fabric_direct_data_i29	: in std_logic := '0';
    fabric_direct_data_i30	: in std_logic := '0';
    fabric_direct_data_i31	: in std_logic := '0';
    fabric_direct_data_i32	: in std_logic := '0';
    fabric_otp_user_pdn_i	: in std_logic := '0';
    fabric_io_oe_i1	: in std_logic := '0';
    fabric_io_oe_i2	: in std_logic := '0';
    fabric_io_oe_i3	: in std_logic := '0';
    fabric_io_oe_i4	: in std_logic := '0';
    fabric_io_oe_i5	: in std_logic := '0';
    fabric_io_oe_i6	: in std_logic := '0';
    fabric_io_oe_i7	: in std_logic := '0';
    fabric_io_oe_i8	: in std_logic := '0';
    fabric_io_oe_i9	: in std_logic := '0';
    fabric_io_oe_i10	: in std_logic := '0';
    fabric_io_oe_i11	: in std_logic := '0';
    fabric_io_oe_i12	: in std_logic := '0';
    fabric_io_oe_i13	: in std_logic := '0';
    fabric_io_oe_i14	: in std_logic := '0';
    fabric_io_oe_i15	: in std_logic := '0';
    fabric_io_oe_i16	: in std_logic := '0';
    fabric_io_oe_i17	: in std_logic := '0';
    fabric_io_oe_i18	: in std_logic := '0';
    fabric_io_oe_i19	: in std_logic := '0';
    fabric_io_oe_i20	: in std_logic := '0';
    fabric_io_oe_i21	: in std_logic := '0';
    fabric_io_oe_i22	: in std_logic := '0';
    fabric_io_oe_i23	: in std_logic := '0';
    fabric_io_oe_i24	: in std_logic := '0';
    fabric_io_oe_i25	: in std_logic := '0';
    fabric_parusr_data_i1	: in std_logic := '0';
    fabric_parusr_data_i2	: in std_logic := '0';
    fabric_parusr_data_i3	: in std_logic := '0';
    fabric_parusr_data_i4	: in std_logic := '0';
    fabric_parusr_data_i5	: in std_logic := '0';
    fabric_parusr_data_i6	: in std_logic := '0';
    fabric_parusr_data_i7	: in std_logic := '0';
    fabric_parusr_data_i8	: in std_logic := '0';
    fabric_parusr_data_i9	: in std_logic := '0';
    fabric_parusr_data_i10	: in std_logic := '0';
    fabric_parusr_data_i11	: in std_logic := '0';
    fabric_parusr_data_i12	: in std_logic := '0';
    fabric_parusr_data_i13	: in std_logic := '0';
    fabric_parusr_data_i14	: in std_logic := '0';
    fabric_parusr_data_i15	: in std_logic := '0';
    fabric_parusr_data_i16	: in std_logic := '0';
    fabric_otp_apb_write_i	: in std_logic := '0';
    fabric_otp_security_testmode_i	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i1	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i2	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i3	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i4	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i5	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i6	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i7	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i8	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i9	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i10	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i11	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i12	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i13	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i14	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i15	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i16	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i17	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i18	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i19	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i20	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i21	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i22	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i23	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i24	: in std_logic := '0';
    fabric_tst_atpg_mrepair_i	: in std_logic := '0';
    fabric_mrepair_fuse_tstscanenable_i	: in std_logic := '0';
    fabric_otp_security_bistmode_i	: in std_logic := '0';
    fabric_lowskew_i22	: in std_logic := '0';
    fabric_lowskew_i23	: in std_logic := '0';
    fabric_lowskew_i20	: in std_logic := '0';
    fabric_otp_user_configreg_i1	: in std_logic := '0';
    fabric_otp_user_configreg_i2	: in std_logic := '0';
    fabric_otp_user_configreg_i3	: in std_logic := '0';
    fabric_otp_user_configreg_i4	: in std_logic := '0';
    fabric_otp_user_configreg_i5	: in std_logic := '0';
    fabric_otp_user_configreg_i6	: in std_logic := '0';
    fabric_otp_user_configreg_i7	: in std_logic := '0';
    fabric_otp_user_configreg_i8	: in std_logic := '0';
    fabric_otp_user_configreg_i9	: in std_logic := '0';
    fabric_otp_user_configreg_i10	: in std_logic := '0';
    fabric_otp_user_configreg_i11	: in std_logic := '0';
    fabric_otp_user_configreg_i12	: in std_logic := '0';
    fabric_otp_user_configreg_i13	: in std_logic := '0';
    fabric_otp_user_configreg_i14	: in std_logic := '0';
    fabric_otp_user_configreg_i15	: in std_logic := '0';
    fabric_otp_user_configreg_i16	: in std_logic := '0';
    fabric_otp_user_configreg_i17	: in std_logic := '0';
    fabric_otp_user_configreg_i18	: in std_logic := '0';
    fabric_otp_user_configreg_i19	: in std_logic := '0';
    fabric_otp_user_configreg_i20	: in std_logic := '0';
    fabric_otp_user_configreg_i21	: in std_logic := '0';
    fabric_otp_user_configreg_i22	: in std_logic := '0';
    fabric_otp_user_configreg_i23	: in std_logic := '0';
    fabric_otp_user_configreg_i24	: in std_logic := '0';
    fabric_otp_user_configreg_i25	: in std_logic := '0';
    fabric_otp_user_configreg_i26	: in std_logic := '0';
    fabric_otp_user_configreg_i27	: in std_logic := '0';
    fabric_otp_user_configreg_i28	: in std_logic := '0';
    fabric_otp_user_configreg_i29	: in std_logic := '0';
    fabric_otp_user_configreg_i30	: in std_logic := '0';
    fabric_otp_user_configreg_i31	: in std_logic := '0';
    fabric_otp_user_configreg_i32	: in std_logic := '0';
    fabric_otp_user_tst_scanin_i1	: in std_logic := '0';
    fabric_otp_user_tst_scanin_i2	: in std_logic := '0';
    fabric_otp_user_tst_scanin_i3	: in std_logic := '0';
    fabric_otp_user_tst_scanin_i4	: in std_logic := '0';
    fabric_otp_user_tst_scanin_i5	: in std_logic := '0';
    fabric_sif_update_en_i1	: in std_logic := '0';
    fabric_sif_update_en_i2	: in std_logic := '0';
    fabric_sif_update_en_i3	: in std_logic := '0';
    fabric_sif_update_en_i4	: in std_logic := '0';
    fabric_sif_update_en_i5	: in std_logic := '0';
    fabric_sif_update_en_i6	: in std_logic := '0';
    fabric_sif_update_en_i7	: in std_logic := '0';
    fabric_sif_update_en_i8	: in std_logic := '0';
    fabric_sif_update_en_i9	: in std_logic := '0';
    fabric_sif_update_en_i10	: in std_logic := '0';
    fabric_sif_update_en_i11	: in std_logic := '0';
    fabric_sif_update_en_i12	: in std_logic := '0';
    fabric_sif_update_en_i13	: in std_logic := '0';
    fabric_sif_update_en_i14	: in std_logic := '0';
    fabric_sif_update_en_i15	: in std_logic := '0';
    fabric_sif_update_en_i16	: in std_logic := '0';
    fabric_sif_update_en_i17	: in std_logic := '0';
    fabric_sif_update_en_i18	: in std_logic := '0';
    fabric_sif_update_en_i19	: in std_logic := '0';
    fabric_sif_update_en_i20	: in std_logic := '0';
    fabric_sif_update_en_i21	: in std_logic := '0';
    fabric_sif_update_en_i22	: in std_logic := '0';
    fabric_sif_update_en_i23	: in std_logic := '0';
    fabric_sif_update_en_i24	: in std_logic := '0';
    fabric_mrepair_por_i	: in std_logic := '0';
    fabric_mrepair_rst_n_i	: in std_logic := '0';
    fabric_mrepair_initn_i	: in std_logic := '0';
    fabric_spare_i1	: in std_logic := '0';
    fabric_spare_i2	: in std_logic := '0';
    fabric_spare_i3	: in std_logic := '0';

    fabric_mrepair_fuse_bbad_o	: out std_logic := '0';
    fabric_jtag_trst_n_o	: out std_logic := '0';
    fabric_debug_direct_permission_write_o1	: out std_logic := '0';
    fabric_debug_direct_permission_write_o2	: out std_logic := '0';
    fabric_debug_direct_permission_write_o3	: out std_logic := '0';
    fabric_debug_direct_permission_write_o4	: out std_logic := '0';
    fabric_otp_security_bist_end1_o	: out std_logic := '0';
    fabric_parusr_data_val_o	: out std_logic := '0';
    fabric_debug_lock_reg_o	: out std_logic := '0';
    fabric_debug_security_error_read_o	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o1	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o2	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o3	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o4	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o5	: out std_logic := '0';
    fabric_otp_user_tst_scanout_o1	: out std_logic := '0';
    fabric_otp_user_tst_scanout_o2	: out std_logic := '0';
    fabric_otp_user_tst_scanout_o3	: out std_logic := '0';
    fabric_otp_user_tst_scanout_o4	: out std_logic := '0';
    fabric_otp_user_tst_scanout_o5	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o1	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o2	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o3	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o4	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o5	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o6	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o7	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o8	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o9	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o10	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o11	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o12	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o13	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o14	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o15	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o16	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o17	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o18	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o19	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o20	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o21	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o22	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o23	: out std_logic := '0';
    fabric_sif_update_en_to_bist_o24	: out std_logic := '0';
    fabric_otp_user_locked_o	: out std_logic := '0';
    fabric_otp_security_bist_bad_o	: out std_logic := '0';
    fabric_debug_frame_permission_frame_o1	: out std_logic := '0';
    fabric_debug_frame_permission_frame_o2	: out std_logic := '0';
    fabric_debug_frame_permission_frame_o3	: out std_logic := '0';
    fabric_debug_frame_permission_frame_o4	: out std_logic := '0';
    fabric_otp_user_pwok_o	: out std_logic := '0';
    fabric_otp_user_bend2_o	: out std_logic := '0';
    fabric_mrepair_fuse_ded_o	: out std_logic := '0';
    fabric_debug_access_reg_data_ready_o	: out std_logic := '0';
    fabric_data_to_bist_o1	: out std_logic := '0';
    fabric_data_to_bist_o2	: out std_logic := '0';
    fabric_data_to_bist_o3	: out std_logic := '0';
    fabric_data_to_bist_o4	: out std_logic := '0';
    fabric_data_to_bist_o5	: out std_logic := '0';
    fabric_data_to_bist_o6	: out std_logic := '0';
    fabric_data_to_bist_o7	: out std_logic := '0';
    fabric_data_to_bist_o8	: out std_logic := '0';
    fabric_data_to_bist_o9	: out std_logic := '0';
    fabric_data_to_bist_o10	: out std_logic := '0';
    fabric_data_to_bist_o11	: out std_logic := '0';
    fabric_data_to_bist_o12	: out std_logic := '0';
    fabric_data_to_bist_o13	: out std_logic := '0';
    fabric_data_to_bist_o14	: out std_logic := '0';
    fabric_data_to_bist_o15	: out std_logic := '0';
    fabric_data_to_bist_o16	: out std_logic := '0';
    fabric_data_to_bist_o17	: out std_logic := '0';
    fabric_data_to_bist_o18	: out std_logic := '0';
    fabric_data_to_bist_o19	: out std_logic := '0';
    fabric_data_to_bist_o20	: out std_logic := '0';
    fabric_data_to_bist_o21	: out std_logic := '0';
    fabric_data_to_bist_o22	: out std_logic := '0';
    fabric_data_to_bist_o23	: out std_logic := '0';
    fabric_data_to_bist_o24	: out std_logic := '0';
    fabric_otp_user_startword_o1	: out std_logic := '0';
    fabric_otp_user_startword_o2	: out std_logic := '0';
    fabric_otp_user_startword_o3	: out std_logic := '0';
    fabric_otp_user_startword_o4	: out std_logic := '0';
    fabric_otp_user_startword_o5	: out std_logic := '0';
    fabric_otp_user_startword_o6	: out std_logic := '0';
    fabric_otp_user_startword_o7	: out std_logic := '0';
    fabric_otp_user_startword_o8	: out std_logic := '0';
    fabric_otp_user_startword_o9	: out std_logic := '0';
    fabric_otp_user_startword_o10	: out std_logic := '0';
    fabric_otp_user_startword_o11	: out std_logic := '0';
    fabric_otp_user_startword_o12	: out std_logic := '0';
    fabric_otp_user_startword_o13	: out std_logic := '0';
    fabric_otp_user_startword_o14	: out std_logic := '0';
    fabric_otp_user_startword_o15	: out std_logic := '0';
    fabric_otp_user_startword_o16	: out std_logic := '0';
    fabric_ahb_direct_data_o1	: out std_logic := '0';
    fabric_ahb_direct_data_o2	: out std_logic := '0';
    fabric_ahb_direct_data_o3	: out std_logic := '0';
    fabric_ahb_direct_data_o4	: out std_logic := '0';
    fabric_ahb_direct_data_o5	: out std_logic := '0';
    fabric_ahb_direct_data_o6	: out std_logic := '0';
    fabric_ahb_direct_data_o7	: out std_logic := '0';
    fabric_ahb_direct_data_o8	: out std_logic := '0';
    fabric_ahb_direct_data_o9	: out std_logic := '0';
    fabric_ahb_direct_data_o10	: out std_logic := '0';
    fabric_ahb_direct_data_o11	: out std_logic := '0';
    fabric_ahb_direct_data_o12	: out std_logic := '0';
    fabric_ahb_direct_data_o13	: out std_logic := '0';
    fabric_ahb_direct_data_o14	: out std_logic := '0';
    fabric_ahb_direct_data_o15	: out std_logic := '0';
    fabric_ahb_direct_data_o16	: out std_logic := '0';
    fabric_ahb_direct_data_o17	: out std_logic := '0';
    fabric_ahb_direct_data_o18	: out std_logic := '0';
    fabric_ahb_direct_data_o19	: out std_logic := '0';
    fabric_ahb_direct_data_o20	: out std_logic := '0';
    fabric_ahb_direct_data_o21	: out std_logic := '0';
    fabric_ahb_direct_data_o22	: out std_logic := '0';
    fabric_ahb_direct_data_o23	: out std_logic := '0';
    fabric_ahb_direct_data_o24	: out std_logic := '0';
    fabric_ahb_direct_data_o25	: out std_logic := '0';
    fabric_ahb_direct_data_o26	: out std_logic := '0';
    fabric_ahb_direct_data_o27	: out std_logic := '0';
    fabric_ahb_direct_data_o28	: out std_logic := '0';
    fabric_ahb_direct_data_o29	: out std_logic := '0';
    fabric_ahb_direct_data_o30	: out std_logic := '0';
    fabric_ahb_direct_data_o31	: out std_logic := '0';
    fabric_ahb_direct_data_o32	: out std_logic := '0';
    fabric_parusr_data_o1	: out std_logic := '0';
    fabric_parusr_data_o2	: out std_logic := '0';
    fabric_parusr_data_o3	: out std_logic := '0';
    fabric_parusr_data_o4	: out std_logic := '0';
    fabric_parusr_data_o5	: out std_logic := '0';
    fabric_parusr_data_o6	: out std_logic := '0';
    fabric_parusr_data_o7	: out std_logic := '0';
    fabric_parusr_data_o8	: out std_logic := '0';
    fabric_parusr_data_o9	: out std_logic := '0';
    fabric_parusr_data_o10	: out std_logic := '0';
    fabric_parusr_data_o11	: out std_logic := '0';
    fabric_parusr_data_o12	: out std_logic := '0';
    fabric_parusr_data_o13	: out std_logic := '0';
    fabric_parusr_data_o14	: out std_logic := '0';
    fabric_parusr_data_o15	: out std_logic := '0';
    fabric_parusr_data_o16	: out std_logic := '0';
    fabric_debug_otp_reload_err_o	: out std_logic := '0';
    fabric_cfg_fabric_user_unmask_o	: out std_logic := '0';
    fabric_decoder_init_ready_o	: out std_logic := '0';
    fabric_global_chip_status_o1	: out std_logic := '0';
    fabric_global_chip_status_o2	: out std_logic := '0';
    fabric_global_chip_status_o3	: out std_logic := '0';
    fabric_debug_security_boot_done_o	: out std_logic := '0';
    fabric_otp_user_calibrated_o	: out std_logic := '0';
    fabric_fuse_status_o1	: out std_logic := '0';
    fabric_fuse_status_o2	: out std_logic := '0';
    fabric_fuse_status_o3	: out std_logic := '0';
    fabric_otp_apb_rdata_o1	: out std_logic := '0';
    fabric_otp_apb_rdata_o2	: out std_logic := '0';
    fabric_otp_apb_rdata_o3	: out std_logic := '0';
    fabric_otp_apb_rdata_o4	: out std_logic := '0';
    fabric_otp_apb_rdata_o5	: out std_logic := '0';
    fabric_otp_apb_rdata_o6	: out std_logic := '0';
    fabric_otp_apb_rdata_o7	: out std_logic := '0';
    fabric_otp_apb_rdata_o8	: out std_logic := '0';
    fabric_otp_apb_rdata_o9	: out std_logic := '0';
    fabric_otp_apb_rdata_o10	: out std_logic := '0';
    fabric_otp_apb_rdata_o11	: out std_logic := '0';
    fabric_otp_apb_rdata_o12	: out std_logic := '0';
    fabric_otp_apb_rdata_o13	: out std_logic := '0';
    fabric_otp_apb_rdata_o14	: out std_logic := '0';
    fabric_otp_apb_rdata_o15	: out std_logic := '0';
    fabric_otp_apb_rdata_o16	: out std_logic := '0';
    fabric_otp_apb_rdata_o17	: out std_logic := '0';
    fabric_otp_apb_rdata_o18	: out std_logic := '0';
    fabric_otp_apb_rdata_o19	: out std_logic := '0';
    fabric_otp_apb_rdata_o20	: out std_logic := '0';
    fabric_otp_apb_rdata_o21	: out std_logic := '0';
    fabric_otp_apb_rdata_o22	: out std_logic := '0';
    fabric_otp_apb_rdata_o23	: out std_logic := '0';
    fabric_otp_apb_rdata_o24	: out std_logic := '0';
    fabric_otp_apb_rdata_o25	: out std_logic := '0';
    fabric_otp_apb_rdata_o26	: out std_logic := '0';
    fabric_otp_apb_rdata_o27	: out std_logic := '0';
    fabric_otp_apb_rdata_o28	: out std_logic := '0';
    fabric_otp_apb_rdata_o29	: out std_logic := '0';
    fabric_otp_apb_rdata_o30	: out std_logic := '0';
    fabric_otp_apb_rdata_o31	: out std_logic := '0';
    fabric_otp_apb_rdata_o32	: out std_logic := '0';
    fabric_jtag_tms_o	: out std_logic := '0';
    fabric_debug_bsec_core_status_o1	: out std_logic := '0';
    fabric_debug_bsec_core_status_o2	: out std_logic := '0';
    fabric_debug_bsec_core_status_o3	: out std_logic := '0';
    fabric_debug_bsec_core_status_o4	: out std_logic := '0';
    fabric_debug_bsec_core_status_o5	: out std_logic := '0';
    fabric_debug_bsec_core_status_o6	: out std_logic := '0';
    fabric_debug_bsec_core_status_o7	: out std_logic := '0';
    fabric_debug_bsec_core_status_o8	: out std_logic := '0';
    fabric_debug_bsec_core_status_o9	: out std_logic := '0';
    fabric_debug_bsec_core_status_o10	: out std_logic := '0';
    fabric_debug_bsec_core_status_o11	: out std_logic := '0';
    fabric_debug_bsec_core_status_o12	: out std_logic := '0';
    fabric_debug_bsec_core_status_o13	: out std_logic := '0';
    fabric_debug_bsec_core_status_o14	: out std_logic := '0';
    fabric_debug_bsec_core_status_o15	: out std_logic := '0';
    fabric_debug_bsec_core_status_o16	: out std_logic := '0';
    fabric_debug_bsec_core_status_o17	: out std_logic := '0';
    fabric_debug_bsec_core_status_o18	: out std_logic := '0';
    fabric_debug_bsec_core_status_o19	: out std_logic := '0';
    fabric_debug_bsec_core_status_o20	: out std_logic := '0';
    fabric_debug_bsec_core_status_o21	: out std_logic := '0';
    fabric_debug_bsec_core_status_o22	: out std_logic := '0';
    fabric_debug_bsec_core_status_o23	: out std_logic := '0';
    fabric_debug_bsec_core_status_o24	: out std_logic := '0';
    fabric_debug_bsec_core_status_o25	: out std_logic := '0';
    fabric_debug_bsec_core_status_o26	: out std_logic := '0';
    fabric_debug_bsec_core_status_o27	: out std_logic := '0';
    fabric_debug_bsec_core_status_o28	: out std_logic := '0';
    fabric_debug_bsec_core_status_o29	: out std_logic := '0';
    fabric_debug_bsec_core_status_o30	: out std_logic := '0';
    fabric_debug_bsec_core_status_o31	: out std_logic := '0';
    fabric_debug_bsec_core_status_o32	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o1	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o2	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o3	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o4	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o5	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o6	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o7	: out std_logic := '0';
    fabric_mrepair_fuse_bist1fail_o8	: out std_logic := '0';
    fabric_flag_ready_o	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o1	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o2	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o3	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o4	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o5	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o6	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o7	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o8	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o9	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o10	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o11	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o12	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o13	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o14	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o15	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o16	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o17	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o18	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o19	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o20	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o21	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o22	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o23	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o24	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o25	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o26	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o27	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o28	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o29	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o30	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o31	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o32	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o33	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o34	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o35	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o36	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o37	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o38	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o39	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o40	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o41	: out std_logic := '0';
    fabric_debug_rst_soft_o	: out std_logic := '0';
    fabric_otp_user_ack_o	: out std_logic := '0';
    fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o	: out std_logic := '0';
    fabric_shift_en_to_bist_o1	: out std_logic := '0';
    fabric_shift_en_to_bist_o2	: out std_logic := '0';
    fabric_shift_en_to_bist_o3	: out std_logic := '0';
    fabric_shift_en_to_bist_o4	: out std_logic := '0';
    fabric_shift_en_to_bist_o5	: out std_logic := '0';
    fabric_shift_en_to_bist_o6	: out std_logic := '0';
    fabric_shift_en_to_bist_o7	: out std_logic := '0';
    fabric_shift_en_to_bist_o8	: out std_logic := '0';
    fabric_shift_en_to_bist_o9	: out std_logic := '0';
    fabric_shift_en_to_bist_o10	: out std_logic := '0';
    fabric_shift_en_to_bist_o11	: out std_logic := '0';
    fabric_shift_en_to_bist_o12	: out std_logic := '0';
    fabric_shift_en_to_bist_o13	: out std_logic := '0';
    fabric_shift_en_to_bist_o14	: out std_logic := '0';
    fabric_shift_en_to_bist_o15	: out std_logic := '0';
    fabric_shift_en_to_bist_o16	: out std_logic := '0';
    fabric_shift_en_to_bist_o17	: out std_logic := '0';
    fabric_shift_en_to_bist_o18	: out std_logic := '0';
    fabric_shift_en_to_bist_o19	: out std_logic := '0';
    fabric_shift_en_to_bist_o20	: out std_logic := '0';
    fabric_shift_en_to_bist_o21	: out std_logic := '0';
    fabric_shift_en_to_bist_o22	: out std_logic := '0';
    fabric_shift_en_to_bist_o23	: out std_logic := '0';
    fabric_shift_en_to_bist_o24	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o1	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o2	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o3	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o4	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o5	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o6	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o7	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o8	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o9	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o10	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o11	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o12	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o13	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o14	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o15	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o16	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o17	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o18	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o19	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o20	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o21	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o22	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o23	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o24	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o25	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o26	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o27	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o28	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o29	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o30	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o31	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o32	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o33	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o34	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o35	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o36	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o37	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o38	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o39	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o40	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o41	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o42	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o43	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o44	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o45	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o46	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o47	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o48	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o49	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o50	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o51	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o52	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o53	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o54	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o55	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o56	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o57	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o58	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o59	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o60	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o61	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o62	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o63	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o64	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o65	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o66	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o67	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o68	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o69	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o70	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o71	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o72	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o73	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o74	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o75	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o76	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o77	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o78	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o79	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o80	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o81	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o82	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o83	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o84	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o85	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o86	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o87	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o88	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o89	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o90	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o91	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o92	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o93	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o94	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o95	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o96	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o97	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o98	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o99	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o100	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o101	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o102	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o103	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o104	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o105	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o106	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o107	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o108	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o109	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o110	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o111	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o112	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o113	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o114	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o115	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o116	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o117	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o118	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o119	: out std_logic := '0';
    fabric_sif_reg_en_to_bist_o120	: out std_logic := '0';
    fabric_debug_otp_manager_read_otp_o	: out std_logic := '0';
    fabric_otp_user_sec_o	: out std_logic := '0';
    fabric_otp_user_wlromout_o1	: out std_logic := '0';
    fabric_otp_user_wlromout_o2	: out std_logic := '0';
    fabric_otp_user_wlromout_o3	: out std_logic := '0';
    fabric_otp_user_wlromout_o4	: out std_logic := '0';
    fabric_otp_user_wlromout_o5	: out std_logic := '0';
    fabric_otp_user_wlromout_o6	: out std_logic := '0';
    fabric_otp_user_wlromout_o7	: out std_logic := '0';
    fabric_otp_user_wlromout_o8	: out std_logic := '0';
    fabric_otp_user_wlromout_o9	: out std_logic := '0';
    fabric_otp_user_wlromout_o10	: out std_logic := '0';
    fabric_mrepair_fuse_bend1_o	: out std_logic := '0';
    fabric_mrepair_fuse_flagstate_o1	: out std_logic := '0';
    fabric_mrepair_fuse_flagstate_o2	: out std_logic := '0';
    fabric_mrepair_fuse_flagstate_o3	: out std_logic := '0';
    fabric_mrepair_fuse_flagstate_o4	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o1	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o2	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o3	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o4	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o5	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o6	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o7	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o8	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o9	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o10	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o11	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o12	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o13	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o14	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o15	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o16	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o17	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o18	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o19	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o20	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o21	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o22	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o23	: out std_logic := '0';
    fabric_system_data_from_mem_bist_o24	: out std_logic := '0';
    fabric_direct_data_o1	: out std_logic := '0';
    fabric_direct_data_o2	: out std_logic := '0';
    fabric_direct_data_o3	: out std_logic := '0';
    fabric_direct_data_o4	: out std_logic := '0';
    fabric_direct_data_o5	: out std_logic := '0';
    fabric_direct_data_o6	: out std_logic := '0';
    fabric_direct_data_o7	: out std_logic := '0';
    fabric_direct_data_o8	: out std_logic := '0';
    fabric_direct_data_o9	: out std_logic := '0';
    fabric_direct_data_o10	: out std_logic := '0';
    fabric_direct_data_o11	: out std_logic := '0';
    fabric_direct_data_o12	: out std_logic := '0';
    fabric_direct_data_o13	: out std_logic := '0';
    fabric_direct_data_o14	: out std_logic := '0';
    fabric_direct_data_o15	: out std_logic := '0';
    fabric_direct_data_o16	: out std_logic := '0';
    fabric_direct_data_o17	: out std_logic := '0';
    fabric_direct_data_o18	: out std_logic := '0';
    fabric_direct_data_o19	: out std_logic := '0';
    fabric_direct_data_o20	: out std_logic := '0';
    fabric_direct_data_o21	: out std_logic := '0';
    fabric_direct_data_o22	: out std_logic := '0';
    fabric_direct_data_o23	: out std_logic := '0';
    fabric_direct_data_o24	: out std_logic := '0';
    fabric_direct_data_o25	: out std_logic := '0';
    fabric_direct_data_o26	: out std_logic := '0';
    fabric_direct_data_o27	: out std_logic := '0';
    fabric_direct_data_o28	: out std_logic := '0';
    fabric_direct_data_o29	: out std_logic := '0';
    fabric_direct_data_o30	: out std_logic := '0';
    fabric_direct_data_o31	: out std_logic := '0';
    fabric_direct_data_o32	: out std_logic := '0';
    fabric_otp_user_bbad_o	: out std_logic := '0';
    fabric_user_read_cycle_o	: out std_logic := '0';
    fabric_chip_status_o1	: out std_logic := '0';
    fabric_chip_status_o2	: out std_logic := '0';
    fabric_chip_status_o3	: out std_logic := '0';
    fabric_chip_status_o4	: out std_logic := '0';
    fabric_chip_status_o5	: out std_logic := '0';
    fabric_chip_status_o6	: out std_logic := '0';
    fabric_chip_status_o7	: out std_logic := '0';
    fabric_chip_status_o8	: out std_logic := '0';
    fabric_chip_status_o9	: out std_logic := '0';
    fabric_chip_status_o10	: out std_logic := '0';
    fabric_chip_status_o11	: out std_logic := '0';
    fabric_chip_status_o12	: out std_logic := '0';
    fabric_chip_status_o13	: out std_logic := '0';
    fabric_chip_status_o14	: out std_logic := '0';
    fabric_chip_status_o15	: out std_logic := '0';
    fabric_chip_status_o16	: out std_logic := '0';
    fabric_chip_status_o17	: out std_logic := '0';
    fabric_chip_status_o18	: out std_logic := '0';
    fabric_chip_status_o19	: out std_logic := '0';
    fabric_chip_status_o20	: out std_logic := '0';
    fabric_chip_status_o21	: out std_logic := '0';
    fabric_chip_status_o22	: out std_logic := '0';
    fabric_chip_status_o23	: out std_logic := '0';
    fabric_chip_status_o24	: out std_logic := '0';
    fabric_chip_status_o25	: out std_logic := '0';
    fabric_chip_status_o26	: out std_logic := '0';
    fabric_chip_status_o27	: out std_logic := '0';
    fabric_chip_status_o28	: out std_logic := '0';
    fabric_chip_status_o29	: out std_logic := '0';
    fabric_chip_status_o30	: out std_logic := '0';
    fabric_chip_status_o31	: out std_logic := '0';
    fabric_chip_status_o32	: out std_logic := '0';
    fabric_chip_status_o33	: out std_logic := '0';
    fabric_chip_status_o34	: out std_logic := '0';
    fabric_chip_status_o35	: out std_logic := '0';
    fabric_chip_status_o36	: out std_logic := '0';
    fabric_chip_status_o37	: out std_logic := '0';
    fabric_chip_status_o38	: out std_logic := '0';
    fabric_chip_status_o39	: out std_logic := '0';
    fabric_chip_status_o40	: out std_logic := '0';
    fabric_chip_status_o41	: out std_logic := '0';
    fabric_chip_status_o42	: out std_logic := '0';
    fabric_chip_status_o43	: out std_logic := '0';
    fabric_chip_status_o44	: out std_logic := '0';
    fabric_chip_status_o45	: out std_logic := '0';
    fabric_chip_status_o46	: out std_logic := '0';
    fabric_chip_status_o47	: out std_logic := '0';
    fabric_chip_status_o48	: out std_logic := '0';
    fabric_chip_status_o49	: out std_logic := '0';
    fabric_chip_status_o50	: out std_logic := '0';
    fabric_chip_status_o51	: out std_logic := '0';
    fabric_chip_status_o52	: out std_logic := '0';
    fabric_chip_status_o53	: out std_logic := '0';
    fabric_chip_status_o54	: out std_logic := '0';
    fabric_chip_status_o55	: out std_logic := '0';
    fabric_chip_status_o56	: out std_logic := '0';
    fabric_chip_status_o57	: out std_logic := '0';
    fabric_chip_status_o58	: out std_logic := '0';
    fabric_chip_status_o59	: out std_logic := '0';
    fabric_chip_status_o60	: out std_logic := '0';
    fabric_chip_status_o61	: out std_logic := '0';
    fabric_chip_status_o62	: out std_logic := '0';
    fabric_chip_status_o63	: out std_logic := '0';
    fabric_chip_status_o64	: out std_logic := '0';
    fabric_chip_status_o65	: out std_logic := '0';
    fabric_chip_status_o66	: out std_logic := '0';
    fabric_chip_status_o67	: out std_logic := '0';
    fabric_chip_status_o68	: out std_logic := '0';
    fabric_chip_status_o69	: out std_logic := '0';
    fabric_chip_status_o70	: out std_logic := '0';
    fabric_chip_status_o71	: out std_logic := '0';
    fabric_chip_status_o72	: out std_logic := '0';
    fabric_mrepair_fuse_disturbed_o	: out std_logic := '0';
    fabric_debug_otpboot_state_o1	: out std_logic := '0';
    fabric_debug_otpboot_state_o2	: out std_logic := '0';
    fabric_debug_otpboot_state_o3	: out std_logic := '0';
    fabric_pd_ready_o1	: out std_logic := '0';
    fabric_pd_ready_o2	: out std_logic := '0';
    fabric_pd_ready_o3	: out std_logic := '0';
    fabric_pd_ready_o4	: out std_logic := '0';
    fabric_pd_ready_o5	: out std_logic := '0';
    fabric_pd_ready_o6	: out std_logic := '0';
    fabric_pd_ready_o7	: out std_logic := '0';
    fabric_pd_ready_o8	: out std_logic := '0';
    fabric_pd_ready_o9	: out std_logic := '0';
    fabric_pd_ready_o10	: out std_logic := '0';
    fabric_pd_ready_o11	: out std_logic := '0';
    fabric_pd_ready_o12	: out std_logic := '0';
    fabric_pd_ready_o13	: out std_logic := '0';
    fabric_pd_ready_o14	: out std_logic := '0';
    fabric_pd_ready_o15	: out std_logic := '0';
    fabric_pd_ready_o16	: out std_logic := '0';
    fabric_pd_ready_o17	: out std_logic := '0';
    fabric_pd_ready_o18	: out std_logic := '0';
    fabric_pd_ready_o19	: out std_logic := '0';
    fabric_pd_ready_o20	: out std_logic := '0';
    fabric_pd_ready_o21	: out std_logic := '0';
    fabric_pd_ready_o22	: out std_logic := '0';
    fabric_pd_ready_o23	: out std_logic := '0';
    fabric_pd_ready_o24	: out std_logic := '0';
    fabric_debug_key_correct_o	: out std_logic := '0';
    fabric_otp_apb_ready_o	: out std_logic := '0';
    fabric_otp_user_progfail_o	: out std_logic := '0';
    fabric_mrepair_fuse_sec_o	: out std_logic := '0';
    fabric_mrepair_fuse_bend2_o	: out std_logic := '0';
    fabric_debug_lifecycle_o1	: out std_logic := '0';
    fabric_debug_lifecycle_o2	: out std_logic := '0';
    fabric_debug_lifecycle_o3	: out std_logic := '0';
    fabric_debug_lifecycle_o4	: out std_logic := '0';
    fabric_mrepair_fuse_ack_o	: out std_logic := '0';
    fabric_debug_cpt_retry_o1	: out std_logic := '0';
    fabric_debug_cpt_retry_o2	: out std_logic := '0';
    fabric_debug_cpt_retry_o3	: out std_logic := '0';
    fabric_debug_cpt_retry_o4	: out std_logic := '0';
    fabric_otp_security_ack_o	: out std_logic := '0';
    fabric_debug_otpmgmt_state_o1	: out std_logic := '0';
    fabric_debug_otpmgmt_state_o2	: out std_logic := '0';
    fabric_debug_otpmgmt_state_o3	: out std_logic := '0';
    fabric_mrepair_fuse_progfail_o	: out std_logic := '0';
    fabric_otp_user_bist2fail_o1	: out std_logic := '0';
    fabric_otp_user_bist2fail_o2	: out std_logic := '0';
    fabric_otp_user_bist2fail_o3	: out std_logic := '0';
    fabric_otp_user_bist2fail_o4	: out std_logic := '0';
    fabric_otp_user_bist2fail_o5	: out std_logic := '0';
    fabric_otp_user_bist2fail_o6	: out std_logic := '0';
    fabric_otp_user_bist2fail_o7	: out std_logic := '0';
    fabric_user_data_o1	: out std_logic := '0';
    fabric_user_data_o2	: out std_logic := '0';
    fabric_user_data_o3	: out std_logic := '0';
    fabric_user_data_o4	: out std_logic := '0';
    fabric_user_data_o5	: out std_logic := '0';
    fabric_user_data_o6	: out std_logic := '0';
    fabric_user_data_o7	: out std_logic := '0';
    fabric_user_data_o8	: out std_logic := '0';
    fabric_user_data_o9	: out std_logic := '0';
    fabric_user_data_o10	: out std_logic := '0';
    fabric_user_data_o11	: out std_logic := '0';
    fabric_user_data_o12	: out std_logic := '0';
    fabric_user_data_o13	: out std_logic := '0';
    fabric_user_data_o14	: out std_logic := '0';
    fabric_user_data_o15	: out std_logic := '0';
    fabric_user_data_o16	: out std_logic := '0';
    fabric_user_data_o17	: out std_logic := '0';
    fabric_user_data_o18	: out std_logic := '0';
    fabric_user_data_o19	: out std_logic := '0';
    fabric_user_data_o20	: out std_logic := '0';
    fabric_user_data_o21	: out std_logic := '0';
    fabric_user_data_o22	: out std_logic := '0';
    fabric_user_data_o23	: out std_logic := '0';
    fabric_user_data_o24	: out std_logic := '0';
    fabric_user_data_o25	: out std_logic := '0';
    fabric_user_data_o26	: out std_logic := '0';
    fabric_user_data_o27	: out std_logic := '0';
    fabric_user_data_o28	: out std_logic := '0';
    fabric_user_data_o29	: out std_logic := '0';
    fabric_user_data_o30	: out std_logic := '0';
    fabric_user_data_o31	: out std_logic := '0';
    fabric_user_data_o32	: out std_logic := '0';
    fabric_jtag_tdi_o	: out std_logic := '0';
    fabric_lowskew_o3	: out std_logic := '0';
    fabric_lowskew_o5	: out std_logic := '0';
    fabric_lowskew_o4	: out std_logic := '0';
    fabric_debug_error_o	: out std_logic := '0';
    fabric_jtag_usr2_o	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o1	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o2	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o3	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o4	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o5	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o6	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o7	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o8	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o9	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o10	: out std_logic := '0';
    fabric_debug_otpapb_state_o1	: out std_logic := '0';
    fabric_debug_otpapb_state_o2	: out std_logic := '0';
    fabric_debug_otpapb_state_o3	: out std_logic := '0';
    fabric_otp_user_bist1fail_o1	: out std_logic := '0';
    fabric_otp_user_bist1fail_o2	: out std_logic := '0';
    fabric_otp_user_bist1fail_o3	: out std_logic := '0';
    fabric_otp_user_bist1fail_o4	: out std_logic := '0';
    fabric_otp_user_bist1fail_o5	: out std_logic := '0';
    fabric_otp_user_bist1fail_o6	: out std_logic := '0';
    fabric_otp_user_bist1fail_o7	: out std_logic := '0';
    fabric_otp_user_bist1fail_o8	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o1	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o2	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o3	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o4	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o5	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o6	: out std_logic := '0';
    fabric_otp_security_bist_fail2_o7	: out std_logic := '0';
    fabric_otp_user_disturbed_o	: out std_logic := '0';
    fabric_flag_trigger_o	: out std_logic := '0';
    fabric_otp_security_bist_end2_o	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o1	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o2	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o3	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o4	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o5	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o6	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o7	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o8	: out std_logic := '0';
    fabric_mrepair_fuse_locked_o	: out std_logic := '0';
    fabric_otp_user_flagstate_o1	: out std_logic := '0';
    fabric_otp_user_flagstate_o2	: out std_logic := '0';
    fabric_otp_user_flagstate_o3	: out std_logic := '0';
    fabric_otp_user_flagstate_o4	: out std_logic := '0';
    fabric_otp_security_scanout_o1	: out std_logic := '0';
    fabric_otp_security_scanout_o2	: out std_logic := '0';
    fabric_otp_security_scanout_o3	: out std_logic := '0';
    fabric_otp_security_scanout_o4	: out std_logic := '0';
    fabric_otp_security_scanout_o5	: out std_logic := '0';
    fabric_user_write_cycle_o	: out std_logic := '0';
    fabric_debug_fsm_state_o1	: out std_logic := '0';
    fabric_debug_fsm_state_o2	: out std_logic := '0';
    fabric_debug_fsm_state_o3	: out std_logic := '0';
    fabric_otp_user_ded_o	: out std_logic := '0';
    fabric_debug_otp_manager_read_done_o	: out std_logic := '0';
    fabric_debug_frame_use_encryption_o	: out std_logic := '0';
    fabric_data_to_system_o	: out std_logic := '0';
    fabric_jtag_usr1_o	: out std_logic := '0';
    fabric_otp_user_bend1_o	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o1	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o2	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o3	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o4	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o5	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o6	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o7	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o8	: out std_logic := '0';
    fabric_mrepair_fuse_ready_o	: out std_logic := '0';
    fabric_mrepair_fuse_calibrated_o	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o1	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o2	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o3	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o4	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o5	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o6	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o7	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o8	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o9	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o10	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o11	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o12	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o13	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o14	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o15	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o16	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o17	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o18	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o19	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o20	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o21	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o22	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o23	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o24	: out std_logic := '0';
    fabric_io_out_o1	: out std_logic := '0';
    fabric_io_out_o2	: out std_logic := '0';
    fabric_io_out_o3	: out std_logic := '0';
    fabric_io_out_o4	: out std_logic := '0';
    fabric_io_out_o5	: out std_logic := '0';
    fabric_io_out_o6	: out std_logic := '0';
    fabric_io_out_o7	: out std_logic := '0';
    fabric_io_out_o8	: out std_logic := '0';
    fabric_io_out_o9	: out std_logic := '0';
    fabric_io_out_o10	: out std_logic := '0';
    fabric_io_out_o11	: out std_logic := '0';
    fabric_io_out_o12	: out std_logic := '0';
    fabric_io_out_o13	: out std_logic := '0';
    fabric_io_out_o14	: out std_logic := '0';
    fabric_io_out_o15	: out std_logic := '0';
    fabric_io_out_o16	: out std_logic := '0';
    fabric_io_out_o17	: out std_logic := '0';
    fabric_io_out_o18	: out std_logic := '0';
    fabric_io_out_o19	: out std_logic := '0';
    fabric_io_out_o20	: out std_logic := '0';
    fabric_io_out_o21	: out std_logic := '0';
    fabric_io_out_o22	: out std_logic := '0';
    fabric_io_out_o23	: out std_logic := '0';
    fabric_io_out_o24	: out std_logic := '0';
    fabric_io_out_o25	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o1	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o2	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o3	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o4	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o5	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o6	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o7	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o8	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o9	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o10	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o11	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o12	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o13	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o14	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o15	: out std_logic := '0';
    fabric_mrepair_fuse_startword_o16	: out std_logic := '0';
    fabric_system_dataready_o	: out std_logic := '0';
    fabric_mrepair_fuse_pwok_o	: out std_logic := '0';
    fabric_lowskew_o6	: out std_logic := '0';
    fabric_cfg_fabric_user_flag_o	: out std_logic := '0';
    fabric_otp_user_dout_o1	: out std_logic := '0';
    fabric_otp_user_dout_o2	: out std_logic := '0';
    fabric_otp_user_dout_o3	: out std_logic := '0';
    fabric_otp_user_dout_o4	: out std_logic := '0';
    fabric_otp_user_dout_o5	: out std_logic := '0';
    fabric_otp_user_dout_o6	: out std_logic := '0';
    fabric_otp_user_dout_o7	: out std_logic := '0';
    fabric_otp_user_dout_o8	: out std_logic := '0';
    fabric_otp_user_dout_o9	: out std_logic := '0';
    fabric_otp_user_dout_o10	: out std_logic := '0';
    fabric_otp_user_dout_o11	: out std_logic := '0';
    fabric_otp_user_dout_o12	: out std_logic := '0';
    fabric_otp_user_dout_o13	: out std_logic := '0';
    fabric_otp_user_dout_o14	: out std_logic := '0';
    fabric_otp_user_dout_o15	: out std_logic := '0';
    fabric_otp_user_dout_o16	: out std_logic := '0';
    fabric_otp_user_dout_o17	: out std_logic := '0';
    fabric_otp_user_dout_o18	: out std_logic := '0';
    fabric_otp_user_dout_o19	: out std_logic := '0';
    fabric_otp_user_dout_o20	: out std_logic := '0';
    fabric_otp_user_dout_o21	: out std_logic := '0';
    fabric_otp_user_dout_o22	: out std_logic := '0';
    fabric_otp_user_dout_o23	: out std_logic := '0';
    fabric_otp_user_dout_o24	: out std_logic := '0';
    fabric_otp_user_dout_o25	: out std_logic := '0';
    fabric_otp_user_dout_o26	: out std_logic := '0';
    fabric_otp_user_dout_o27	: out std_logic := '0';
    fabric_otp_user_dout_o28	: out std_logic := '0';
    fabric_otp_user_dout_o29	: out std_logic := '0';
    fabric_otp_user_dout_o30	: out std_logic := '0';
    fabric_otp_user_dout_o31	: out std_logic := '0';
    fabric_otp_user_dout_o32	: out std_logic := '0';
    fabric_otp_user_dout_o33	: out std_logic := '0';
    fabric_otp_user_dout_o34	: out std_logic := '0';
    fabric_otp_user_dout_o35	: out std_logic := '0';
    fabric_otp_user_dout_o36	: out std_logic := '0';
    fabric_otp_user_dout_o37	: out std_logic := '0';
    fabric_otp_user_dout_o38	: out std_logic := '0';
    fabric_otp_user_dout_o39	: out std_logic := '0';
    fabric_otp_user_dout_o40	: out std_logic := '0';
    fabric_otp_user_dout_o41	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o1	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o2	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o3	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o4	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o5	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o6	: out std_logic := '0';
    fabric_mrepair_fuse_bist2fail_o7	: out std_logic := '0';
    fabric_status_cold_start_o	: out std_logic := '0';
    fabric_flag_error_o	: out std_logic := '0';
    fabric_debug_direct_permission_read_o1	: out std_logic := '0';
    fabric_debug_direct_permission_read_o2	: out std_logic := '0';
    fabric_debug_direct_permission_read_o3	: out std_logic := '0';
    fabric_debug_direct_permission_read_o4	: out std_logic := '0'
);
end component NX_SERVICE_U;

component NX_SERVICE_U_WRAP is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    fabric_otp_user_tst_scanenable_i	: in std_logic := '0';
    fabric_otp_cfg_loader_read_en_i	: in std_logic := '0';
    fabric_otp_security_force_pdn1_i	: in std_logic := '0';
    fabric_otp_security_scanenable_i	: in std_logic := '0';
    fabric_otp_user_din_i	: in std_logic_vector(38 downto 0) := (others => '0');
    fabric_mrepair_fuse_prgwidth_i	: in std_logic_vector(2 downto 0) := (others => '0');
    fabric_otp_apb_wdata_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_cfg_clk_otpm_disable_i	: in std_logic := '0';
    fabric_otp_user_disturbcheck_i	: in std_logic := '0';
    fabric_mrepair_fuse_read_i	: in std_logic := '0';
    fabric_otp_user_rbact2_i	: in std_logic := '0';
    fabric_mrepair_fuse_eccbypass_i	: in std_logic := '0';
    fabric_otp_user_bistmode_i	: in std_logic := '0';
    fabric_otp_user_add_i	: in std_logic_vector(6 downto 0) := (others => '0');
    fabric_otp_user_tm_i	: in std_logic := '0';
    fabric_otp_rstn_i	: in std_logic := '0';
    fabric_mrepair_fuse_disturbchecked_i	: in std_logic := '0';
    fabric_otp_user_rbact1_i	: in std_logic := '0';
    fabric_mrepair_fuse_tst_scanin_i	: in std_logic_vector(4 downto 0) := (others => '0');
    fabric_parusr_type_i	: in std_logic_vector(1 downto 0) := (others => '0');
    fabric_mrepair_fuse_redbypass_i	: in std_logic := '0';
    fabric_otp_user_eccbypass_i	: in std_logic := '0';
    fabric_otp_user_redbypass_i	: in std_logic := '0';
    fabric_mrepair_mode_i	: in std_logic_vector(3 downto 0) := (others => '0');
    fabric_parusr_cs_i	: in std_logic := '0';
    fabric_sif_reg_en_i	: in std_logic_vector(119 downto 0) := (others => '0');
    fabric_mrepair_fuse_rbact2_i	: in std_logic := '0';
    fabric_data_from_system_i	: in std_logic := '0';
    fabric_data_from_bist_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_otp_apb_enable_i	: in std_logic := '0';
    fabric_mrepair_fuse_tm_i	: in std_logic := '0';
    fabric_otp_security_rbact2_i	: in std_logic := '0';
    fabric_otp_security_rbact1_i	: in std_logic := '0';
    fabric_shift_en_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_otp_cfg_loader_write_en_i	: in std_logic := '0';
    fabric_user_data_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_mrepair_fuse_suppadd_i	: in std_logic := '0';
    fabric_mrepair_fuse_prog_i	: in std_logic := '0';
    fabric_otp_user_wordlock_i	: in std_logic := '0';
    fabric_ahb_direct_data_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_user_prog_i	: in std_logic := '0';
    fabric_pd_active_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_otp_user_suppadd_i	: in std_logic := '0';
    fabric_mrepair_fuse_pdn_i	: in std_logic := '0';
    fabric_otp_security_scanin_i	: in std_logic_vector(4 downto 0) := (others => '0');
    fabric_end_encoding_i	: in std_logic := '0';
    fabric_jtag_tdo_usr2_i	: in std_logic := '0';
    fabric_mrepair_fuse_wordlock_i	: in std_logic := '0';
    fabric_otp_user_prgwidth_i	: in std_logic_vector(2 downto 0) := (others => '0');
    fabric_otp_user_read_i	: in std_logic := '0';
    fabric_mrepair_fuse_add_i	: in std_logic_vector(6 downto 0) := (others => '0');
    fabric_mrepair_fuse_bistmode_i	: in std_logic := '0';
    fabric_jtag_tdo_usr1_i	: in std_logic := '0';
    fabric_otp_cfg_clk_fab_en_i	: in std_logic := '0';
    fabric_io_in_i	: in std_logic_vector(24 downto 0) := (others => '0');
    fabric_sif_load_en_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_mrepair_fuse_din_i	: in std_logic_vector(38 downto 0) := (others => '0');
    fabric_otp_apb_addr_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_apb_sel_i	: in std_logic := '0';
    fabric_mrepair_fuse_rbact1_i	: in std_logic := '0';
    fabric_mrepair_fuse_configreg_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_cfg_fabric_apb_en_i	: in std_logic := '0';
    fabric_data_shift_en_i	: in std_logic := '0';
    fabric_lowskew_i21	: in std_logic := '0';
    fabric_direct_data_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_user_pdn_i	: in std_logic := '0';
    fabric_io_oe_i	: in std_logic_vector(24 downto 0) := (others => '0');
    fabric_parusr_data_i	: in std_logic_vector(15 downto 0) := (others => '0');
    fabric_otp_apb_write_i	: in std_logic := '0';
    fabric_otp_security_testmode_i	: in std_logic := '0';
    fabric_system_data_to_mem_bist_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_tst_atpg_mrepair_i	: in std_logic := '0';
    fabric_mrepair_fuse_tstscanenable_i	: in std_logic := '0';
    fabric_otp_security_bistmode_i	: in std_logic := '0';
    fabric_lowskew_i22	: in std_logic := '0';
    fabric_lowskew_i23	: in std_logic := '0';
    fabric_lowskew_i20	: in std_logic := '0';
    fabric_otp_user_configreg_i	: in std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_user_tst_scanin_i	: in std_logic_vector(4 downto 0) := (others => '0');
    fabric_sif_update_en_i	: in std_logic_vector(23 downto 0) := (others => '0');
    fabric_mrepair_por_i	: in std_logic := '0';
    fabric_mrepair_rst_n_i	: in std_logic := '0';
    fabric_mrepair_initn_i	: in std_logic := '0';
    fabric_spare_i	: in std_logic_vector(2 downto 0) := (others => '0');

    fabric_mrepair_fuse_bbad_o	: out std_logic := '0';
    fabric_jtag_trst_n_o	: out std_logic := '0';
    fabric_debug_direct_permission_write_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_otp_security_bist_end1_o	: out std_logic := '0';
    fabric_parusr_data_val_o	: out std_logic := '0';
    fabric_debug_lock_reg_o	: out std_logic := '0';
    fabric_debug_security_error_read_o	: out std_logic := '0';
    fabric_mrepair_fuse_tstscanout_o	: out std_logic_vector(4 downto 0) := (others => '0');
    fabric_otp_user_tst_scanout_o	: out std_logic_vector(4 downto 0) := (others => '0');
    fabric_sif_update_en_to_bist_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_otp_user_locked_o	: out std_logic := '0';
    fabric_otp_security_bist_bad_o	: out std_logic := '0';
    fabric_debug_frame_permission_frame_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_otp_user_pwok_o	: out std_logic := '0';
    fabric_otp_user_bend2_o	: out std_logic := '0';
    fabric_mrepair_fuse_ded_o	: out std_logic := '0';
    fabric_debug_access_reg_data_ready_o	: out std_logic := '0';
    fabric_data_to_bist_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_otp_user_startword_o	: out std_logic_vector(15 downto 0) := (others => '0');
    fabric_ahb_direct_data_o	: out std_logic_vector(31 downto 0) := (others => '0');
    fabric_parusr_data_o	: out std_logic_vector(15 downto 0) := (others => '0');
    fabric_debug_otp_reload_err_o	: out std_logic := '0';
    fabric_cfg_fabric_user_unmask_o	: out std_logic := '0';
    fabric_decoder_init_ready_o	: out std_logic := '0';
    fabric_global_chip_status_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_debug_security_boot_done_o	: out std_logic := '0';
    fabric_otp_user_calibrated_o	: out std_logic := '0';
    fabric_fuse_status_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_otp_apb_rdata_o	: out std_logic_vector(31 downto 0) := (others => '0');
    fabric_jtag_tms_o	: out std_logic := '0';
    fabric_debug_bsec_core_status_o	: out std_logic_vector(31 downto 0) := (others => '0');
    fabric_mrepair_fuse_bist1fail_o	: out std_logic_vector(7 downto 0) := (others => '0');
    fabric_flag_ready_o	: out std_logic := '0';
    fabric_mrepair_fuse_dout_o	: out std_logic_vector(40 downto 0) := (others => '0');
    fabric_debug_rst_soft_o	: out std_logic := '0';
    fabric_otp_user_ack_o	: out std_logic := '0';
    fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o	: out std_logic := '0';
    fabric_shift_en_to_bist_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_sif_reg_en_to_bist_o	: out std_logic_vector(119 downto 0) := (others => '0');
    fabric_debug_otp_manager_read_otp_o	: out std_logic := '0';
    fabric_otp_user_sec_o	: out std_logic := '0';
    fabric_otp_user_wlromout_o	: out std_logic_vector(9 downto 0) := (others => '0');
    fabric_mrepair_fuse_bend1_o	: out std_logic := '0';
    fabric_mrepair_fuse_flagstate_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_system_data_from_mem_bist_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_direct_data_o	: out std_logic_vector(31 downto 0) := (others => '0');
    fabric_otp_user_bbad_o	: out std_logic := '0';
    fabric_user_read_cycle_o	: out std_logic := '0';
    fabric_chip_status_o	: out std_logic_vector(71 downto 0) := (others => '0');
    fabric_mrepair_fuse_disturbed_o	: out std_logic := '0';
    fabric_debug_otpboot_state_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_pd_ready_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_debug_key_correct_o	: out std_logic := '0';
    fabric_otp_apb_ready_o	: out std_logic := '0';
    fabric_otp_user_progfail_o	: out std_logic := '0';
    fabric_mrepair_fuse_sec_o	: out std_logic := '0';
    fabric_mrepair_fuse_bend2_o	: out std_logic := '0';
    fabric_debug_lifecycle_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_mrepair_fuse_ack_o	: out std_logic := '0';
    fabric_debug_cpt_retry_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_otp_security_ack_o	: out std_logic := '0';
    fabric_debug_otpmgmt_state_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_mrepair_fuse_progfail_o	: out std_logic := '0';
    fabric_otp_user_bist2fail_o	: out std_logic_vector(6 downto 0) := (others => '0');
    fabric_user_data_o	: out std_logic_vector(31 downto 0) := (others => '0');
    fabric_jtag_tdi_o	: out std_logic := '0';
    fabric_lowskew_o3	: out std_logic := '0';
    fabric_lowskew_o5	: out std_logic := '0';
    fabric_lowskew_o4	: out std_logic := '0';
    fabric_debug_error_o	: out std_logic := '0';
    fabric_jtag_usr2_o	: out std_logic := '0';
    fabric_mrepair_fuse_wlromout_o	: out std_logic_vector(9 downto 0) := (others => '0');
    fabric_debug_otpapb_state_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_otp_user_bist1fail_o	: out std_logic_vector(7 downto 0) := (others => '0');
    fabric_otp_security_bist_fail2_o	: out std_logic_vector(6 downto 0) := (others => '0');
    fabric_otp_user_disturbed_o	: out std_logic := '0';
    fabric_flag_trigger_o	: out std_logic := '0';
    fabric_otp_security_bist_end2_o	: out std_logic := '0';
    fabric_otp_security_bist_fail1_o	: out std_logic_vector(7 downto 0) := (others => '0');
    fabric_mrepair_fuse_locked_o	: out std_logic := '0';
    fabric_otp_user_flagstate_o	: out std_logic_vector(3 downto 0) := (others => '0');
    fabric_otp_security_scanout_o	: out std_logic_vector(4 downto 0) := (others => '0');
    fabric_user_write_cycle_o	: out std_logic := '0';
    fabric_debug_fsm_state_o	: out std_logic_vector(2 downto 0) := (others => '0');
    fabric_otp_user_ded_o	: out std_logic := '0';
    fabric_debug_otp_manager_read_done_o	: out std_logic := '0';
    fabric_debug_frame_use_encryption_o	: out std_logic := '0';
    fabric_data_to_system_o	: out std_logic := '0';
    fabric_jtag_usr1_o	: out std_logic := '0';
    fabric_otp_user_bend1_o	: out std_logic := '0';
    fabric_debug_otpboot_curr_addr_o	: out std_logic_vector(7 downto 0) := (others => '0');
    fabric_mrepair_fuse_ready_o	: out std_logic := '0';
    fabric_mrepair_fuse_calibrated_o	: out std_logic := '0';
    fabric_sif_load_en_to_bist_o	: out std_logic_vector(23 downto 0) := (others => '0');
    fabric_io_out_o	: out std_logic_vector(24 downto 0) := (others => '0');
    fabric_mrepair_fuse_startword_o	: out std_logic_vector(15 downto 0) := (others => '0');
    fabric_system_dataready_o	: out std_logic := '0';
    fabric_mrepair_fuse_pwok_o	: out std_logic := '0';
    fabric_lowskew_o6	: out std_logic := '0';
    fabric_cfg_fabric_user_flag_o	: out std_logic := '0';
    fabric_otp_user_dout_o	: out std_logic_vector(40 downto 0) := (others => '0');
    fabric_mrepair_fuse_bist2fail_o	: out std_logic_vector(6 downto 0) := (others => '0');
    fabric_status_cold_start_o	: out std_logic := '0';
    fabric_flag_error_o	: out std_logic := '0';
    fabric_debug_direct_permission_read_o	: out std_logic_vector(3 downto 0) := (others => '0')
);
end component NX_SERVICE_U_WRAP;

component NX_SOC_INTERFACE is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    -- dahlia <-> fabric
    fabric_lowskew_o1	: out std_logic := '0';
    fabric_lowskew_i1	: in std_logic := '0';
    fabric_lowskew_i2	: in std_logic := '0';
    fabric_lowskew_i3	: in std_logic := '0';
    fabric_lowskew_i4	: in std_logic := '0';
    fabric_lowskew_i5	: in std_logic := '0';
    fabric_lowskew_i6	: in std_logic := '0';
    fabric_lowskew_i7	: in std_logic := '0';
    fabric_lowskew_i8	: in std_logic := '0';
    fabric_lowskew_i9	: in std_logic := '0';
    fabric_lowskew_i10	: in std_logic := '0';
    fabric_lowskew_o2	: out std_logic := '0';
    fabric_fpga_nic_rstn_i1	: in std_logic := '0';
    fabric_fpga_nic_rstn_i2	: in std_logic := '0';
    fabric_fpga_nic_rstn_i3	: in std_logic := '0';
    fabric_fpga_nic_rstn_i4	: in std_logic := '0';
    fabric_fpga_nic_rstn_i5	: in std_logic := '0';
    fabric_fpga_nic_rstn_i6	: in std_logic := '0';
    fabric_fpga_nic_rstn_i7	: in std_logic := '0';
    fabric_fpga_nic_rstn_i8	: in std_logic := '0';
    fabric_fpga_nic_rstn_i9	: in std_logic := '0';
    fabric_fpga_nic_rstn_i10	: in std_logic := '0';
    fabric_fpga_pmrstn_i	: in std_logic := '0';
    fabric_fpga_sysrstn_i	: in std_logic := '0';
    fabric_fpga_trigger_in_o1	: out std_logic := '0';
    fabric_fpga_trigger_in_o2	: out std_logic := '0';
    fabric_fpga_trigger_in_o3	: out std_logic := '0';
    fabric_fpga_trigger_in_o4	: out std_logic := '0';
    fabric_fpga_trigger_in_o5	: out std_logic := '0';
    fabric_fpga_trigger_in_o6	: out std_logic := '0';
    fabric_fpga_trigger_in_o7	: out std_logic := '0';
    fabric_fpga_trigger_in_o8	: out std_logic := '0';
    fabric_fpga_trigger_out_i1	: in std_logic := '0';
    fabric_fpga_trigger_out_i2	: in std_logic := '0';
    fabric_fpga_trigger_out_i3	: in std_logic := '0';
    fabric_fpga_trigger_out_i4	: in std_logic := '0';
    fabric_fpga_trigger_out_i5	: in std_logic := '0';
    fabric_fpga_trigger_out_i6	: in std_logic := '0';
    fabric_fpga_trigger_out_i7	: in std_logic := '0';
    fabric_fpga_trigger_out_i8	: in std_logic := '0';
    fabric_fpga_interrupt_in_i1	: in std_logic := '0';
    fabric_fpga_interrupt_in_i2	: in std_logic := '0';
    fabric_fpga_interrupt_in_i3	: in std_logic := '0';
    fabric_fpga_interrupt_in_i4	: in std_logic := '0';
    fabric_fpga_interrupt_in_i5	: in std_logic := '0';
    fabric_fpga_interrupt_in_i6	: in std_logic := '0';
    fabric_fpga_interrupt_in_i7	: in std_logic := '0';
    fabric_fpga_interrupt_in_i8	: in std_logic := '0';
    fabric_fpga_interrupt_in_i9	: in std_logic := '0';
    fabric_fpga_interrupt_in_i10	: in std_logic := '0';
    fabric_fpga_interrupt_in_i11	: in std_logic := '0';
    fabric_fpga_interrupt_in_i12	: in std_logic := '0';
    fabric_fpga_interrupt_in_i13	: in std_logic := '0';
    fabric_fpga_interrupt_in_i14	: in std_logic := '0';
    fabric_fpga_interrupt_in_i15	: in std_logic := '0';
    fabric_fpga_interrupt_in_i16	: in std_logic := '0';
    fabric_fpga_interrupt_in_i17	: in std_logic := '0';
    fabric_fpga_interrupt_in_i18	: in std_logic := '0';
    fabric_fpga_interrupt_in_i19	: in std_logic := '0';
    fabric_fpga_interrupt_in_i20	: in std_logic := '0';
    fabric_fpga_interrupt_in_i21	: in std_logic := '0';
    fabric_fpga_interrupt_in_i22	: in std_logic := '0';
    fabric_fpga_interrupt_in_i23	: in std_logic := '0';
    fabric_fpga_interrupt_in_i24	: in std_logic := '0';
    fabric_fpga_interrupt_in_i25	: in std_logic := '0';
    fabric_fpga_interrupt_in_i26	: in std_logic := '0';
    fabric_fpga_interrupt_in_i27	: in std_logic := '0';
    fabric_fpga_interrupt_in_i28	: in std_logic := '0';
    fabric_fpga_interrupt_in_i29	: in std_logic := '0';
    fabric_fpga_interrupt_in_i30	: in std_logic := '0';
    fabric_fpga_interrupt_in_i31	: in std_logic := '0';
    fabric_fpga_interrupt_in_i32	: in std_logic := '0';
    fabric_fpga_interrupt_in_i33	: in std_logic := '0';
    fabric_fpga_interrupt_in_i34	: in std_logic := '0';
    fabric_fpga_interrupt_in_i35	: in std_logic := '0';
    fabric_fpga_interrupt_in_i36	: in std_logic := '0';
    fabric_fpga_interrupt_in_i37	: in std_logic := '0';
    fabric_fpga_interrupt_in_i38	: in std_logic := '0';
    fabric_fpga_interrupt_in_i39	: in std_logic := '0';
    fabric_fpga_interrupt_in_i40	: in std_logic := '0';
    fabric_fpga_interrupt_in_i41	: in std_logic := '0';
    fabric_fpga_interrupt_in_i42	: in std_logic := '0';
    fabric_fpga_interrupt_in_i43	: in std_logic := '0';
    fabric_fpga_interrupt_in_i44	: in std_logic := '0';
    fabric_fpga_interrupt_in_i45	: in std_logic := '0';
    fabric_fpga_interrupt_in_i46	: in std_logic := '0';
    fabric_fpga_interrupt_in_i47	: in std_logic := '0';
    fabric_fpga_interrupt_in_i48	: in std_logic := '0';
    fabric_fpga_interrupt_in_i49	: in std_logic := '0';
    fabric_fpga_interrupt_in_i50	: in std_logic := '0';
    fabric_fpga_interrupt_in_i51	: in std_logic := '0';
    fabric_fpga_interrupt_in_i52	: in std_logic := '0';
    fabric_fpga_interrupt_in_i53	: in std_logic := '0';
    fabric_fpga_interrupt_in_i54	: in std_logic := '0';
    fabric_fpga_interrupt_in_i55	: in std_logic := '0';
    fabric_fpga_interrupt_in_i56	: in std_logic := '0';
    fabric_fpga_interrupt_in_i57	: in std_logic := '0';
    fabric_fpga_interrupt_in_i58	: in std_logic := '0';
    fabric_fpga_interrupt_in_i59	: in std_logic := '0';
    fabric_fpga_interrupt_in_i60	: in std_logic := '0';
    fabric_fpga_interrupt_in_i61	: in std_logic := '0';
    fabric_fpga_interrupt_in_i62	: in std_logic := '0';
    fabric_fpga_interrupt_in_i63	: in std_logic := '0';
    fabric_fpga_interrupt_in_i64	: in std_logic := '0';
    fabric_fpga_interrupt_in_i65	: in std_logic := '0';
    fabric_fpga_interrupt_in_i66	: in std_logic := '0';
    fabric_fpga_interrupt_in_i67	: in std_logic := '0';
    fabric_fpga_interrupt_in_i68	: in std_logic := '0';
    fabric_fpga_interrupt_in_i69	: in std_logic := '0';
    fabric_fpga_interrupt_in_i70	: in std_logic := '0';
    fabric_fpga_interrupt_in_i71	: in std_logic := '0';
    fabric_fpga_interrupt_in_i72	: in std_logic := '0';
    fabric_fpga_interrupt_in_i73	: in std_logic := '0';
    fabric_fpga_interrupt_in_i74	: in std_logic := '0';
    fabric_fpga_interrupt_in_i75	: in std_logic := '0';
    fabric_fpga_interrupt_in_i76	: in std_logic := '0';
    fabric_fpga_interrupt_in_i77	: in std_logic := '0';
    fabric_fpga_interrupt_in_i78	: in std_logic := '0';
    fabric_fpga_interrupt_in_i79	: in std_logic := '0';
    fabric_fpga_interrupt_in_i80	: in std_logic := '0';
    fabric_fpga_interrupt_in_i81	: in std_logic := '0';
    fabric_fpga_interrupt_in_i82	: in std_logic := '0';
    fabric_fpga_interrupt_in_i83	: in std_logic := '0';
    fabric_fpga_interrupt_in_i84	: in std_logic := '0';
    fabric_fpga_interrupt_in_i85	: in std_logic := '0';
    fabric_fpga_interrupt_in_i86	: in std_logic := '0';
    fabric_fpga_interrupt_in_i87	: in std_logic := '0';
    fabric_fpga_interrupt_in_i88	: in std_logic := '0';
    fabric_fpga_interrupt_in_i89	: in std_logic := '0';
    fabric_fpga_interrupt_in_i90	: in std_logic := '0';
    fabric_fpga_interrupt_in_i91	: in std_logic := '0';
    fabric_fpga_interrupt_in_i92	: in std_logic := '0';
    fabric_fpga_interrupt_in_i93	: in std_logic := '0';
    fabric_fpga_interrupt_in_i94	: in std_logic := '0';
    fabric_fpga_interrupt_in_i95	: in std_logic := '0';
    fabric_fpga_interrupt_in_i96	: in std_logic := '0';
    fabric_fpga_interrupt_in_i97	: in std_logic := '0';
    fabric_fpga_interrupt_in_i98	: in std_logic := '0';
    fabric_fpga_interrupt_in_i99	: in std_logic := '0';
    fabric_fpga_interrupt_in_i100	: in std_logic := '0';
    fabric_fpga_interrupt_in_i101	: in std_logic := '0';
    fabric_fpga_interrupt_in_i102	: in std_logic := '0';
    fabric_fpga_interrupt_in_i103	: in std_logic := '0';
    fabric_fpga_interrupt_in_i104	: in std_logic := '0';
    fabric_fpga_interrupt_in_i105	: in std_logic := '0';
    fabric_fpga_interrupt_in_i106	: in std_logic := '0';
    fabric_fpga_interrupt_in_i107	: in std_logic := '0';
    fabric_fpga_interrupt_in_i108	: in std_logic := '0';
    fabric_fpga_interrupt_in_i109	: in std_logic := '0';
    fabric_fpga_interrupt_in_i110	: in std_logic := '0';
    fabric_fpga_interrupt_in_i111	: in std_logic := '0';
    fabric_fpga_interrupt_in_i112	: in std_logic := '0';
    fabric_fpga_interrupt_in_i113	: in std_logic := '0';
    fabric_fpga_interrupt_in_i114	: in std_logic := '0';
    fabric_fpga_interrupt_in_i115	: in std_logic := '0';
    fabric_fpga_interrupt_in_i116	: in std_logic := '0';
    fabric_fpga_interrupt_in_i117	: in std_logic := '0';
    fabric_fpga_interrupt_in_i118	: in std_logic := '0';
    fabric_fpga_interrupt_in_i119	: in std_logic := '0';
    fabric_fpga_interrupt_in_i120	: in std_logic := '0';
    fabric_sysc_hold_on_debug_i	: in std_logic := '0';
    fabric_fpga_events60_i1	: in std_logic := '0';
    fabric_fpga_events60_i2	: in std_logic := '0';
    fabric_fpga_events60_i3	: in std_logic := '0';
    fabric_fpga_events60_i4	: in std_logic := '0';
    fabric_fpga_events60_i5	: in std_logic := '0';
    fabric_fpga_events60_i6	: in std_logic := '0';
    fabric_fpga_events60_i7	: in std_logic := '0';
    fabric_fpga_events60_i8	: in std_logic := '0';
    fabric_fpga_events60_i9	: in std_logic := '0';
    fabric_fpga_events60_i10	: in std_logic := '0';
    fabric_fpga_events60_i11	: in std_logic := '0';
    fabric_fpga_events60_i12	: in std_logic := '0';
    fabric_fpga_events60_i13	: in std_logic := '0';
    fabric_fpga_events60_i14	: in std_logic := '0';
    fabric_fpga_events60_i15	: in std_logic := '0';
    fabric_fpga_events60_i16	: in std_logic := '0';
    fabric_fpga_events60_i17	: in std_logic := '0';
    fabric_fpga_events60_i18	: in std_logic := '0';
    fabric_fpga_events60_i19	: in std_logic := '0';
    fabric_fpga_events60_i20	: in std_logic := '0';
    fabric_fpga_events60_i21	: in std_logic := '0';
    fabric_fpga_events60_i22	: in std_logic := '0';
    fabric_fpga_events60_i23	: in std_logic := '0';
    fabric_fpga_events60_i24	: in std_logic := '0';
    fabric_fpga_events60_i25	: in std_logic := '0';
    fabric_fpga_events60_i26	: in std_logic := '0';
    fabric_fpga_events60_i27	: in std_logic := '0';
    fabric_fpga_events60_i28	: in std_logic := '0';
    fabric_fpga_events60_i29	: in std_logic := '0';
    fabric_fpga_events60_i30	: in std_logic := '0';
    fabric_fpga_events60_i31	: in std_logic := '0';
    fabric_fpga_events60_i32	: in std_logic := '0';
    fabric_fpga_events60_i33	: in std_logic := '0';
    fabric_fpga_events60_i34	: in std_logic := '0';
    fabric_fpga_events60_i35	: in std_logic := '0';
    fabric_fpga_events60_i36	: in std_logic := '0';
    fabric_fpga_events60_i37	: in std_logic := '0';
    fabric_fpga_events60_i38	: in std_logic := '0';
    fabric_fpga_events60_i39	: in std_logic := '0';
    fabric_fpga_events60_i40	: in std_logic := '0';
    fabric_fpga_events60_i41	: in std_logic := '0';
    fabric_fpga_events60_i42	: in std_logic := '0';
    fabric_fpga_events60_i43	: in std_logic := '0';
    fabric_fpga_events60_i44	: in std_logic := '0';
    fabric_fpga_events60_i45	: in std_logic := '0';
    fabric_fpga_events60_i46	: in std_logic := '0';
    fabric_fpga_events60_i47	: in std_logic := '0';
    fabric_fpga_events60_i48	: in std_logic := '0';
    fabric_fpga_events60_i49	: in std_logic := '0';
    fabric_fpga_events60_i50	: in std_logic := '0';
    fabric_fpga_events60_i51	: in std_logic := '0';
    fabric_fpga_events60_i52	: in std_logic := '0';
    fabric_fpga_events60_i53	: in std_logic := '0';
    fabric_fpga_events60_i54	: in std_logic := '0';
    fabric_fpga_events60_i55	: in std_logic := '0';
    fabric_fpga_events60_i56	: in std_logic := '0';
    fabric_fpga_events60_i57	: in std_logic := '0';
    fabric_fpga_events60_i58	: in std_logic := '0';
    fabric_fpga_events60_i59	: in std_logic := '0';
    fabric_fpga_events60_i60	: in std_logic := '0';
    fabric_fpga_araddr_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o13	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o14	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o15	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o16	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o17	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o18	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o19	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o20	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o21	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o22	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o23	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o24	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o25	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o26	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o27	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o28	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o29	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o30	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o31	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o32	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o33	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o34	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o35	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o36	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o37	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o38	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o39	: out std_logic := '0';
    fabric_fpga_araddr_axi_s1_o40	: out std_logic := '0';
    fabric_fpga_arburst_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arburst_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arcache_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arcache_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arcache_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arcache_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_arid_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_arlen_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_arlock_axi_s1_o	: out std_logic := '0';
    fabric_fpga_arprot_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arprot_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arprot_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arqos_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arqos_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arqos_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arqos_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_arregion_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arregion_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arregion_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arregion_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_arsize_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_arsize_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_arsize_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_arvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o13	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o14	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o15	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o16	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o17	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o18	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o19	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o20	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o21	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o22	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o23	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o24	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o25	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o26	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o27	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o28	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o29	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o30	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o31	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o32	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o33	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o34	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o35	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o36	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o37	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o38	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o39	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o40	: out std_logic := '0';
    fabric_fpga_awburst_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awburst_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awcache_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awcache_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awcache_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awcache_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_awid_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_awlen_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_awlock_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awprot_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awprot_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awprot_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awqos_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awqos_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awqos_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awqos_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awregion_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awregion_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awregion_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_awregion_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_awsize_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_awsize_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_awsize_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_bready_axi_s1_o	: out std_logic := '0';
    fabric_fpga_rready_axi_s1_o	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o13	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o14	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o15	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o16	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o17	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o18	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o19	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o20	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o21	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o22	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o23	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o24	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o25	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o26	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o27	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o28	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o29	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o30	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o31	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o32	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o33	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o34	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o35	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o36	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o37	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o38	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o39	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o40	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o41	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o42	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o43	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o44	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o45	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o46	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o47	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o48	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o49	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o50	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o51	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o52	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o53	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o54	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o55	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o56	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o57	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o58	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o59	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o60	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o61	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o62	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o63	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o64	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o65	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o66	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o67	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o68	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o69	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o70	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o71	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o72	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o73	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o74	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o75	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o76	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o77	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o78	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o79	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o80	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o81	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o82	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o83	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o84	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o85	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o86	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o87	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o88	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o89	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o90	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o91	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o92	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o93	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o94	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o95	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o96	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o97	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o98	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o99	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o100	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o101	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o102	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o103	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o104	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o105	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o106	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o107	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o108	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o109	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o110	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o111	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o112	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o113	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o114	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o115	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o116	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o117	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o118	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o119	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o120	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o121	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o122	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o123	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o124	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o125	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o126	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o127	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o128	: out std_logic := '0';
    fabric_fpga_wlast_axi_s1_o	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o1	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o2	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o3	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o4	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o5	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o6	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o7	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o8	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o9	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o10	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o11	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o12	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o13	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o14	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o15	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o16	: out std_logic := '0';
    fabric_fpga_wvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_arready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_awready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i1	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i2	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i3	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i4	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i5	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i6	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i7	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i8	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i9	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i10	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i11	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i12	: in std_logic := '0';
    fabric_fpga_bresp_axi_s1_i1	: in std_logic := '0';
    fabric_fpga_bresp_axi_s1_i2	: in std_logic := '0';
    fabric_fpga_bvalid_axi_s1_i	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i1	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i2	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i3	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i4	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i5	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i6	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i7	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i8	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i9	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i10	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i11	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i12	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i13	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i14	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i15	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i16	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i17	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i18	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i19	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i20	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i21	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i22	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i23	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i24	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i25	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i26	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i27	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i28	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i29	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i30	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i31	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i32	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i33	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i34	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i35	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i36	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i37	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i38	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i39	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i40	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i41	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i42	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i43	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i44	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i45	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i46	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i47	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i48	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i49	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i50	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i51	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i52	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i53	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i54	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i55	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i56	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i57	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i58	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i59	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i60	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i61	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i62	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i63	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i64	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i65	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i66	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i67	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i68	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i69	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i70	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i71	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i72	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i73	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i74	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i75	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i76	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i77	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i78	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i79	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i80	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i81	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i82	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i83	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i84	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i85	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i86	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i87	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i88	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i89	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i90	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i91	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i92	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i93	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i94	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i95	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i96	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i97	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i98	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i99	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i100	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i101	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i102	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i103	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i104	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i105	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i106	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i107	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i108	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i109	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i110	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i111	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i112	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i113	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i114	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i115	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i116	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i117	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i118	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i119	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i120	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i121	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i122	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i123	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i124	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i125	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i126	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i127	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i128	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i1	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i2	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i3	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i4	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i5	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i6	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i7	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i8	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i9	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i10	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i11	: in std_logic := '0';
    fabric_fpga_rid_axi_s1_i12	: in std_logic := '0';
    fabric_fpga_rlast_axi_s1_i	: in std_logic := '0';
    fabric_fpga_rresp_axi_s1_i1	: in std_logic := '0';
    fabric_fpga_rresp_axi_s1_i2	: in std_logic := '0';
    fabric_fpga_rvalid_axi_s1_i	: in std_logic := '0';
    fabric_fpga_wready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_araddr_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o13	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o14	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o15	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o16	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o17	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o18	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o19	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o20	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o21	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o22	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o23	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o24	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o25	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o26	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o27	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o28	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o29	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o30	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o31	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o32	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o33	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o34	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o35	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o36	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o37	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o38	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o39	: out std_logic := '0';
    fabric_fpga_araddr_axi_s2_o40	: out std_logic := '0';
    fabric_fpga_arburst_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arburst_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arcache_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arcache_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arcache_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arcache_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_arid_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_arlen_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_arlock_axi_s2_o	: out std_logic := '0';
    fabric_fpga_arprot_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arprot_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arprot_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arqos_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arqos_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arqos_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arqos_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_arregion_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arregion_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arregion_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arregion_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_arsize_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_arsize_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_arsize_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_arvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o13	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o14	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o15	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o16	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o17	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o18	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o19	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o20	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o21	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o22	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o23	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o24	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o25	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o26	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o27	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o28	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o29	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o30	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o31	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o32	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o33	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o34	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o35	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o36	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o37	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o38	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o39	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o40	: out std_logic := '0';
    fabric_fpga_awburst_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awburst_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awcache_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awcache_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awcache_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awcache_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_awid_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_awlen_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_awlock_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awprot_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awprot_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awprot_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awqos_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awqos_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awqos_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awqos_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awregion_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awregion_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awregion_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_awregion_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_awsize_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_awsize_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_awsize_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_bready_axi_s2_o	: out std_logic := '0';
    fabric_fpga_rready_axi_s2_o	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o13	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o14	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o15	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o16	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o17	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o18	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o19	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o20	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o21	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o22	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o23	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o24	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o25	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o26	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o27	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o28	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o29	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o30	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o31	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o32	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o33	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o34	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o35	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o36	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o37	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o38	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o39	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o40	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o41	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o42	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o43	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o44	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o45	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o46	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o47	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o48	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o49	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o50	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o51	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o52	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o53	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o54	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o55	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o56	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o57	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o58	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o59	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o60	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o61	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o62	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o63	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o64	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o65	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o66	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o67	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o68	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o69	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o70	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o71	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o72	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o73	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o74	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o75	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o76	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o77	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o78	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o79	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o80	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o81	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o82	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o83	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o84	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o85	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o86	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o87	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o88	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o89	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o90	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o91	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o92	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o93	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o94	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o95	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o96	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o97	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o98	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o99	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o100	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o101	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o102	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o103	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o104	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o105	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o106	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o107	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o108	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o109	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o110	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o111	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o112	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o113	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o114	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o115	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o116	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o117	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o118	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o119	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o120	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o121	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o122	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o123	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o124	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o125	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o126	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o127	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o128	: out std_logic := '0';
    fabric_fpga_wlast_axi_s2_o	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o1	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o2	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o3	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o4	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o5	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o6	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o7	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o8	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o9	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o10	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o11	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o12	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o13	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o14	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o15	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o16	: out std_logic := '0';
    fabric_fpga_wvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_arready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_awready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i1	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i2	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i3	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i4	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i5	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i6	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i7	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i8	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i9	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i10	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i11	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i12	: in std_logic := '0';
    fabric_fpga_bresp_axi_s2_i1	: in std_logic := '0';
    fabric_fpga_bresp_axi_s2_i2	: in std_logic := '0';
    fabric_fpga_bvalid_axi_s2_i	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i1	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i2	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i3	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i4	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i5	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i6	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i7	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i8	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i9	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i10	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i11	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i12	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i13	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i14	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i15	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i16	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i17	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i18	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i19	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i20	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i21	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i22	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i23	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i24	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i25	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i26	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i27	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i28	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i29	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i30	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i31	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i32	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i33	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i34	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i35	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i36	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i37	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i38	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i39	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i40	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i41	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i42	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i43	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i44	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i45	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i46	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i47	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i48	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i49	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i50	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i51	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i52	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i53	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i54	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i55	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i56	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i57	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i58	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i59	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i60	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i61	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i62	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i63	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i64	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i65	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i66	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i67	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i68	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i69	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i70	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i71	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i72	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i73	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i74	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i75	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i76	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i77	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i78	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i79	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i80	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i81	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i82	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i83	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i84	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i85	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i86	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i87	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i88	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i89	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i90	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i91	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i92	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i93	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i94	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i95	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i96	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i97	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i98	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i99	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i100	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i101	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i102	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i103	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i104	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i105	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i106	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i107	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i108	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i109	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i110	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i111	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i112	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i113	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i114	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i115	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i116	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i117	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i118	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i119	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i120	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i121	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i122	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i123	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i124	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i125	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i126	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i127	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i128	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i1	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i2	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i3	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i4	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i5	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i6	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i7	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i8	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i9	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i10	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i11	: in std_logic := '0';
    fabric_fpga_rid_axi_s2_i12	: in std_logic := '0';
    fabric_fpga_rlast_axi_s2_i	: in std_logic := '0';
    fabric_fpga_rresp_axi_s2_i1	: in std_logic := '0';
    fabric_fpga_rresp_axi_s2_i2	: in std_logic := '0';
    fabric_fpga_rvalid_axi_s2_i	: in std_logic := '0';
    fabric_fpga_wready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_arready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_awready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o1	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o2	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o3	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o4	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o5	: out std_logic := '0';
    fabric_fpga_bresp_axi_m1_o1	: out std_logic := '0';
    fabric_fpga_bresp_axi_m1_o2	: out std_logic := '0';
    fabric_fpga_bvalid_axi_m1_o	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o1	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o2	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o3	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o4	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o5	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o6	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o1	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o2	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o3	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o4	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o5	: out std_logic := '0';
    fabric_fpga_dma_finish_m1_o6	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o1	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o2	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o3	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o4	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o5	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o6	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o7	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o8	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o9	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o10	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o11	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o12	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o13	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o14	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o15	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o16	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o17	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o18	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o19	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o20	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o21	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o22	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o23	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o24	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o25	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o26	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o27	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o28	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o29	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o30	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o31	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o32	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o33	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o34	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o35	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o36	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o37	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o38	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o39	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o40	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o41	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o42	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o43	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o44	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o45	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o46	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o47	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o48	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o49	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o50	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o51	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o52	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o53	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o54	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o55	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o56	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o57	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o58	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o59	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o60	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o61	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o62	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o63	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o64	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o65	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o66	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o67	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o68	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o69	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o70	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o71	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o72	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o73	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o74	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o75	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o76	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o77	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o78	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o79	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o80	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o81	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o82	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o83	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o84	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o85	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o86	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o87	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o88	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o89	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o90	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o91	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o92	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o93	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o94	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o95	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o96	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o97	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o98	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o99	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o100	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o101	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o102	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o103	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o104	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o105	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o106	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o107	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o108	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o109	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o110	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o111	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o112	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o113	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o114	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o115	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o116	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o117	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o118	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o119	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o120	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o121	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o122	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o123	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o124	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o125	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o126	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o127	: out std_logic := '0';
    fabric_fpga_rdata_axi_m1_o128	: out std_logic := '0';
    fabric_fpga_rid_axi_m1_o1	: out std_logic := '0';
    fabric_fpga_rid_axi_m1_o2	: out std_logic := '0';
    fabric_fpga_rid_axi_m1_o3	: out std_logic := '0';
    fabric_fpga_rid_axi_m1_o4	: out std_logic := '0';
    fabric_fpga_rid_axi_m1_o5	: out std_logic := '0';
    fabric_fpga_rlast_axi_m1_o	: out std_logic := '0';
    fabric_fpga_rresp_axi_m1_o1	: out std_logic := '0';
    fabric_fpga_rresp_axi_m1_o2	: out std_logic := '0';
    fabric_fpga_rvalid_axi_m1_o	: out std_logic := '0';
    fabric_fpga_wready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_araddr_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i9	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i10	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i11	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i12	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i13	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i14	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i15	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i16	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i17	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i18	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i19	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i20	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i21	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i22	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i23	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i24	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i25	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i26	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i27	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i28	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i29	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i30	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i31	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i32	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i33	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i34	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i35	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i36	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i37	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i38	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i39	: in std_logic := '0';
    fabric_fpga_araddr_axi_m1_i40	: in std_logic := '0';
    fabric_fpga_arburst_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arburst_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arcache_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arcache_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arcache_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arcache_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_arid_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arid_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arid_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arid_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_arid_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_arlen_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_arlock_axi_m1_i	: in std_logic := '0';
    fabric_fpga_arprot_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arprot_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arprot_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arqos_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arqos_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arqos_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arqos_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_arsize_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_arsize_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_arsize_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_arvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i9	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i10	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i11	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i12	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i13	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i14	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i15	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i16	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i17	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i18	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i19	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i20	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i21	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i22	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i23	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i24	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i25	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i26	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i27	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i28	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i29	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i30	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i31	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i32	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i33	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i34	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i35	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i36	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i37	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i38	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i39	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i40	: in std_logic := '0';
    fabric_fpga_awburst_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awburst_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awcache_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awcache_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awcache_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awcache_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_awid_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awid_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awid_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awid_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_awid_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_awlen_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_awlock_axi_m1_i	: in std_logic := '0';
    fabric_fpga_awprot_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awprot_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awprot_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awqos_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awqos_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awqos_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awqos_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_awsize_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_awsize_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_awsize_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_awvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_bready_axi_m1_i	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i1	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i2	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i3	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i4	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i5	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i6	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i1	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i2	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i3	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i4	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i5	: in std_logic := '0';
    fabric_fpga_dma_req_m1_i6	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i1	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i2	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i3	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i4	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i5	: in std_logic := '0';
    fabric_fpga_dma_single_m1_i6	: in std_logic := '0';
    fabric_fpga_rready_axi_m1_i	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i9	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i10	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i11	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i12	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i13	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i14	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i15	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i16	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i17	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i18	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i19	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i20	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i21	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i22	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i23	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i24	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i25	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i26	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i27	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i28	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i29	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i30	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i31	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i32	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i33	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i34	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i35	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i36	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i37	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i38	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i39	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i40	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i41	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i42	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i43	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i44	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i45	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i46	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i47	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i48	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i49	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i50	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i51	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i52	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i53	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i54	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i55	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i56	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i57	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i58	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i59	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i60	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i61	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i62	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i63	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i64	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i65	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i66	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i67	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i68	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i69	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i70	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i71	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i72	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i73	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i74	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i75	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i76	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i77	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i78	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i79	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i80	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i81	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i82	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i83	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i84	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i85	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i86	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i87	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i88	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i89	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i90	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i91	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i92	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i93	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i94	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i95	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i96	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i97	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i98	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i99	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i100	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i101	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i102	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i103	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i104	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i105	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i106	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i107	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i108	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i109	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i110	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i111	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i112	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i113	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i114	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i115	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i116	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i117	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i118	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i119	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i120	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i121	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i122	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i123	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i124	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i125	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i126	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i127	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i128	: in std_logic := '0';
    fabric_fpga_wlast_axi_m1_i	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i1	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i2	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i3	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i4	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i5	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i6	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i7	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i8	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i9	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i10	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i11	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i12	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i13	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i14	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i15	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i16	: in std_logic := '0';
    fabric_fpga_wvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_arready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_awready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o1	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o2	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o3	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o4	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o5	: out std_logic := '0';
    fabric_fpga_bresp_axi_m2_o1	: out std_logic := '0';
    fabric_fpga_bresp_axi_m2_o2	: out std_logic := '0';
    fabric_fpga_bvalid_axi_m2_o	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o1	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o2	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o3	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o4	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o5	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o6	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o1	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o2	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o3	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o4	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o5	: out std_logic := '0';
    fabric_fpga_dma_finish_m2_o6	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o1	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o2	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o3	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o4	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o5	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o6	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o7	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o8	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o9	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o10	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o11	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o12	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o13	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o14	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o15	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o16	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o17	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o18	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o19	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o20	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o21	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o22	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o23	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o24	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o25	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o26	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o27	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o28	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o29	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o30	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o31	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o32	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o33	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o34	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o35	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o36	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o37	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o38	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o39	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o40	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o41	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o42	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o43	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o44	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o45	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o46	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o47	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o48	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o49	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o50	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o51	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o52	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o53	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o54	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o55	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o56	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o57	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o58	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o59	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o60	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o61	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o62	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o63	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o64	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o65	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o66	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o67	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o68	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o69	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o70	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o71	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o72	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o73	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o74	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o75	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o76	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o77	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o78	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o79	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o80	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o81	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o82	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o83	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o84	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o85	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o86	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o87	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o88	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o89	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o90	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o91	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o92	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o93	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o94	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o95	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o96	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o97	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o98	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o99	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o100	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o101	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o102	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o103	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o104	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o105	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o106	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o107	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o108	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o109	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o110	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o111	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o112	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o113	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o114	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o115	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o116	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o117	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o118	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o119	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o120	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o121	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o122	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o123	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o124	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o125	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o126	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o127	: out std_logic := '0';
    fabric_fpga_rdata_axi_m2_o128	: out std_logic := '0';
    fabric_fpga_rid_axi_m2_o1	: out std_logic := '0';
    fabric_fpga_rid_axi_m2_o2	: out std_logic := '0';
    fabric_fpga_rid_axi_m2_o3	: out std_logic := '0';
    fabric_fpga_rid_axi_m2_o4	: out std_logic := '0';
    fabric_fpga_rid_axi_m2_o5	: out std_logic := '0';
    fabric_fpga_rlast_axi_m2_o	: out std_logic := '0';
    fabric_fpga_rresp_axi_m2_o1	: out std_logic := '0';
    fabric_fpga_rresp_axi_m2_o2	: out std_logic := '0';
    fabric_fpga_rvalid_axi_m2_o	: out std_logic := '0';
    fabric_fpga_wready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_araddr_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i9	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i10	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i11	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i12	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i13	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i14	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i15	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i16	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i17	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i18	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i19	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i20	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i21	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i22	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i23	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i24	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i25	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i26	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i27	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i28	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i29	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i30	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i31	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i32	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i33	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i34	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i35	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i36	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i37	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i38	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i39	: in std_logic := '0';
    fabric_fpga_araddr_axi_m2_i40	: in std_logic := '0';
    fabric_fpga_arburst_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arburst_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arcache_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arcache_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arcache_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arcache_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_arid_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arid_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arid_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arid_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_arid_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_arlen_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_arlock_axi_m2_i	: in std_logic := '0';
    fabric_fpga_arprot_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arprot_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arprot_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arqos_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arqos_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arqos_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arqos_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_arsize_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_arsize_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_arsize_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_arvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i9	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i10	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i11	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i12	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i13	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i14	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i15	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i16	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i17	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i18	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i19	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i20	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i21	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i22	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i23	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i24	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i25	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i26	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i27	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i28	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i29	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i30	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i31	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i32	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i33	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i34	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i35	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i36	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i37	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i38	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i39	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i40	: in std_logic := '0';
    fabric_fpga_awburst_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awburst_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awcache_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awcache_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awcache_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awcache_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_awid_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awid_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awid_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awid_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_awid_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_awlen_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_awlock_axi_m2_i	: in std_logic := '0';
    fabric_fpga_awprot_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awprot_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awprot_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awqos_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awqos_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awqos_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awqos_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_awsize_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_awsize_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_awsize_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_awvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_bready_axi_m2_i	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i1	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i2	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i3	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i4	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i5	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i6	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i1	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i2	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i3	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i4	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i5	: in std_logic := '0';
    fabric_fpga_dma_req_m2_i6	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i1	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i2	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i3	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i4	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i5	: in std_logic := '0';
    fabric_fpga_dma_single_m2_i6	: in std_logic := '0';
    fabric_fpga_rready_axi_m2_i	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i9	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i10	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i11	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i12	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i13	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i14	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i15	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i16	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i17	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i18	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i19	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i20	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i21	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i22	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i23	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i24	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i25	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i26	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i27	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i28	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i29	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i30	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i31	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i32	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i33	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i34	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i35	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i36	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i37	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i38	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i39	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i40	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i41	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i42	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i43	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i44	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i45	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i46	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i47	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i48	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i49	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i50	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i51	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i52	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i53	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i54	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i55	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i56	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i57	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i58	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i59	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i60	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i61	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i62	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i63	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i64	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i65	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i66	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i67	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i68	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i69	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i70	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i71	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i72	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i73	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i74	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i75	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i76	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i77	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i78	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i79	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i80	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i81	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i82	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i83	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i84	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i85	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i86	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i87	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i88	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i89	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i90	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i91	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i92	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i93	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i94	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i95	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i96	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i97	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i98	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i99	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i100	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i101	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i102	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i103	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i104	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i105	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i106	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i107	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i108	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i109	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i110	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i111	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i112	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i113	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i114	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i115	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i116	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i117	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i118	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i119	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i120	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i121	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i122	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i123	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i124	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i125	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i126	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i127	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i128	: in std_logic := '0';
    fabric_fpga_wlast_axi_m2_i	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i1	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i2	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i3	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i4	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i5	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i6	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i7	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i8	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i9	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i10	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i11	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i12	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i13	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i14	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i15	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i16	: in std_logic := '0';
    fabric_fpga_wvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_ddr0_arready_o	: out std_logic := '0';
    fabric_fpga_ddr0_awready_o	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o1	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o2	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o3	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o4	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o5	: out std_logic := '0';
    fabric_fpga_ddr0_bresp_o1	: out std_logic := '0';
    fabric_fpga_ddr0_bresp_o2	: out std_logic := '0';
    fabric_fpga_ddr0_bvalid_o	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o1	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o2	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o3	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o4	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o5	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o6	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o7	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o8	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o9	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o10	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o11	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o12	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o13	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o14	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o15	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o16	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o17	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o18	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o19	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o20	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o21	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o22	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o23	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o24	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o25	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o26	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o27	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o28	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o29	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o30	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o31	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o32	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o33	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o34	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o35	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o36	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o37	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o38	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o39	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o40	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o41	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o42	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o43	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o44	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o45	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o46	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o47	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o48	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o49	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o50	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o51	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o52	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o53	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o54	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o55	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o56	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o57	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o58	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o59	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o60	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o61	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o62	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o63	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o64	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o65	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o66	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o67	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o68	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o69	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o70	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o71	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o72	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o73	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o74	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o75	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o76	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o77	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o78	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o79	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o80	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o81	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o82	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o83	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o84	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o85	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o86	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o87	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o88	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o89	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o90	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o91	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o92	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o93	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o94	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o95	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o96	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o97	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o98	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o99	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o100	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o101	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o102	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o103	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o104	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o105	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o106	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o107	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o108	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o109	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o110	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o111	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o112	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o113	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o114	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o115	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o116	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o117	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o118	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o119	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o120	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o121	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o122	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o123	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o124	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o125	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o126	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o127	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o128	: out std_logic := '0';
    fabric_fpga_ddr0_rid_o1	: out std_logic := '0';
    fabric_fpga_ddr0_rid_o2	: out std_logic := '0';
    fabric_fpga_ddr0_rid_o3	: out std_logic := '0';
    fabric_fpga_ddr0_rid_o4	: out std_logic := '0';
    fabric_fpga_ddr0_rid_o5	: out std_logic := '0';
    fabric_fpga_ddr0_rlast_o	: out std_logic := '0';
    fabric_fpga_ddr0_rresp_o1	: out std_logic := '0';
    fabric_fpga_ddr0_rresp_o2	: out std_logic := '0';
    fabric_fpga_ddr0_rvalid_o	: out std_logic := '0';
    fabric_fpga_ddr0_wready_o	: out std_logic := '0';
    fabric_fpga_ddr0_araddr_i1	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i2	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i3	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i4	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i5	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i6	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i7	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i8	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i9	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i10	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i11	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i12	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i13	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i14	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i15	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i16	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i17	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i18	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i19	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i20	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i21	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i22	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i23	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i24	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i25	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i26	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i27	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i28	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i29	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i30	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i31	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i32	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i33	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i34	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i35	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i36	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i37	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i38	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i39	: in std_logic := '0';
    fabric_fpga_ddr0_araddr_i40	: in std_logic := '0';
    fabric_fpga_ddr0_arburst_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arburst_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arcache_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arcache_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arcache_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arcache_i4	: in std_logic := '0';
    fabric_fpga_ddr0_arid_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arid_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arid_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arid_i4	: in std_logic := '0';
    fabric_fpga_ddr0_arid_i5	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i4	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i5	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i6	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i7	: in std_logic := '0';
    fabric_fpga_ddr0_arlen_i8	: in std_logic := '0';
    fabric_fpga_ddr0_arlock_i	: in std_logic := '0';
    fabric_fpga_ddr0_arprot_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arprot_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arprot_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arqos_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arqos_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arqos_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arqos_i4	: in std_logic := '0';
    fabric_fpga_ddr0_arsize_i1	: in std_logic := '0';
    fabric_fpga_ddr0_arsize_i2	: in std_logic := '0';
    fabric_fpga_ddr0_arsize_i3	: in std_logic := '0';
    fabric_fpga_ddr0_arvalid_i	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i4	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i5	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i6	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i7	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i8	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i9	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i10	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i11	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i12	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i13	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i14	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i15	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i16	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i17	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i18	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i19	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i20	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i21	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i22	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i23	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i24	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i25	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i26	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i27	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i28	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i29	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i30	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i31	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i32	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i33	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i34	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i35	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i36	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i37	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i38	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i39	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i40	: in std_logic := '0';
    fabric_fpga_ddr0_awburst_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awburst_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awcache_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awcache_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awcache_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awcache_i4	: in std_logic := '0';
    fabric_fpga_ddr0_awid_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awid_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awid_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awid_i4	: in std_logic := '0';
    fabric_fpga_ddr0_awid_i5	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i4	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i5	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i6	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i7	: in std_logic := '0';
    fabric_fpga_ddr0_awlen_i8	: in std_logic := '0';
    fabric_fpga_ddr0_awlock_i	: in std_logic := '0';
    fabric_fpga_ddr0_awprot_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awprot_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awprot_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awqos_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awqos_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awqos_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awqos_i4	: in std_logic := '0';
    fabric_fpga_ddr0_awsize_i1	: in std_logic := '0';
    fabric_fpga_ddr0_awsize_i2	: in std_logic := '0';
    fabric_fpga_ddr0_awsize_i3	: in std_logic := '0';
    fabric_fpga_ddr0_awvalid_i	: in std_logic := '0';
    fabric_fpga_ddr0_bready_i	: in std_logic := '0';
    fabric_fpga_ddr0_rready_i	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i1	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i2	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i3	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i4	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i5	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i6	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i7	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i8	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i9	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i10	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i11	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i12	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i13	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i14	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i15	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i16	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i17	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i18	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i19	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i20	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i21	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i22	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i23	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i24	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i25	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i26	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i27	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i28	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i29	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i30	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i31	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i32	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i33	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i34	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i35	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i36	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i37	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i38	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i39	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i40	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i41	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i42	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i43	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i44	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i45	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i46	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i47	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i48	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i49	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i50	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i51	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i52	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i53	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i54	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i55	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i56	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i57	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i58	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i59	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i60	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i61	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i62	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i63	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i64	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i65	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i66	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i67	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i68	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i69	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i70	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i71	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i72	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i73	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i74	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i75	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i76	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i77	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i78	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i79	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i80	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i81	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i82	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i83	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i84	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i85	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i86	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i87	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i88	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i89	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i90	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i91	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i92	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i93	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i94	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i95	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i96	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i97	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i98	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i99	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i100	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i101	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i102	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i103	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i104	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i105	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i106	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i107	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i108	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i109	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i110	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i111	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i112	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i113	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i114	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i115	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i116	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i117	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i118	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i119	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i120	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i121	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i122	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i123	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i124	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i125	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i126	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i127	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i128	: in std_logic := '0';
    fabric_fpga_ddr0_wlast_i	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i1	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i2	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i3	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i4	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i5	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i6	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i7	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i8	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i9	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i10	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i11	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i12	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i13	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i14	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i15	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i16	: in std_logic := '0';
    fabric_fpga_ddr0_wvalid_i	: in std_logic := '0';
    fabric_fpga_paddr_apb_o1	: out std_logic := '0';
    fabric_fpga_paddr_apb_o2	: out std_logic := '0';
    fabric_fpga_paddr_apb_o3	: out std_logic := '0';
    fabric_fpga_paddr_apb_o4	: out std_logic := '0';
    fabric_fpga_paddr_apb_o5	: out std_logic := '0';
    fabric_fpga_paddr_apb_o6	: out std_logic := '0';
    fabric_fpga_paddr_apb_o7	: out std_logic := '0';
    fabric_fpga_paddr_apb_o8	: out std_logic := '0';
    fabric_fpga_paddr_apb_o9	: out std_logic := '0';
    fabric_fpga_paddr_apb_o10	: out std_logic := '0';
    fabric_fpga_paddr_apb_o11	: out std_logic := '0';
    fabric_fpga_paddr_apb_o12	: out std_logic := '0';
    fabric_fpga_paddr_apb_o13	: out std_logic := '0';
    fabric_fpga_paddr_apb_o14	: out std_logic := '0';
    fabric_fpga_paddr_apb_o15	: out std_logic := '0';
    fabric_fpga_paddr_apb_o16	: out std_logic := '0';
    fabric_fpga_paddr_apb_o17	: out std_logic := '0';
    fabric_fpga_paddr_apb_o18	: out std_logic := '0';
    fabric_fpga_paddr_apb_o19	: out std_logic := '0';
    fabric_fpga_paddr_apb_o20	: out std_logic := '0';
    fabric_fpga_paddr_apb_o21	: out std_logic := '0';
    fabric_fpga_paddr_apb_o22	: out std_logic := '0';
    fabric_fpga_paddr_apb_o23	: out std_logic := '0';
    fabric_fpga_paddr_apb_o24	: out std_logic := '0';
    fabric_fpga_paddr_apb_o25	: out std_logic := '0';
    fabric_fpga_paddr_apb_o26	: out std_logic := '0';
    fabric_fpga_paddr_apb_o27	: out std_logic := '0';
    fabric_fpga_paddr_apb_o28	: out std_logic := '0';
    fabric_fpga_paddr_apb_o29	: out std_logic := '0';
    fabric_fpga_paddr_apb_o30	: out std_logic := '0';
    fabric_fpga_paddr_apb_o31	: out std_logic := '0';
    fabric_fpga_paddr_apb_o32	: out std_logic := '0';
    fabric_fpga_penable_apb_o	: out std_logic := '0';
    fabric_fpga_psel_apb_o	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o1	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o2	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o3	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o4	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o5	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o6	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o7	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o8	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o9	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o10	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o11	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o12	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o13	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o14	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o15	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o16	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o17	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o18	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o19	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o20	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o21	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o22	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o23	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o24	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o25	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o26	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o27	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o28	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o29	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o30	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o31	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o32	: out std_logic := '0';
    fabric_fpga_pwrite_apb_o	: out std_logic := '0';
    fabric_fpga_prdata_apb_i1	: in std_logic := '0';
    fabric_fpga_prdata_apb_i2	: in std_logic := '0';
    fabric_fpga_prdata_apb_i3	: in std_logic := '0';
    fabric_fpga_prdata_apb_i4	: in std_logic := '0';
    fabric_fpga_prdata_apb_i5	: in std_logic := '0';
    fabric_fpga_prdata_apb_i6	: in std_logic := '0';
    fabric_fpga_prdata_apb_i7	: in std_logic := '0';
    fabric_fpga_prdata_apb_i8	: in std_logic := '0';
    fabric_fpga_prdata_apb_i9	: in std_logic := '0';
    fabric_fpga_prdata_apb_i10	: in std_logic := '0';
    fabric_fpga_prdata_apb_i11	: in std_logic := '0';
    fabric_fpga_prdata_apb_i12	: in std_logic := '0';
    fabric_fpga_prdata_apb_i13	: in std_logic := '0';
    fabric_fpga_prdata_apb_i14	: in std_logic := '0';
    fabric_fpga_prdata_apb_i15	: in std_logic := '0';
    fabric_fpga_prdata_apb_i16	: in std_logic := '0';
    fabric_fpga_prdata_apb_i17	: in std_logic := '0';
    fabric_fpga_prdata_apb_i18	: in std_logic := '0';
    fabric_fpga_prdata_apb_i19	: in std_logic := '0';
    fabric_fpga_prdata_apb_i20	: in std_logic := '0';
    fabric_fpga_prdata_apb_i21	: in std_logic := '0';
    fabric_fpga_prdata_apb_i22	: in std_logic := '0';
    fabric_fpga_prdata_apb_i23	: in std_logic := '0';
    fabric_fpga_prdata_apb_i24	: in std_logic := '0';
    fabric_fpga_prdata_apb_i25	: in std_logic := '0';
    fabric_fpga_prdata_apb_i26	: in std_logic := '0';
    fabric_fpga_prdata_apb_i27	: in std_logic := '0';
    fabric_fpga_prdata_apb_i28	: in std_logic := '0';
    fabric_fpga_prdata_apb_i29	: in std_logic := '0';
    fabric_fpga_prdata_apb_i30	: in std_logic := '0';
    fabric_fpga_prdata_apb_i31	: in std_logic := '0';
    fabric_fpga_prdata_apb_i32	: in std_logic := '0';
    fabric_fpga_pready_apb_i	: in std_logic := '0';
    fabric_fpga_pslverr_apb_i	: in std_logic := '0';
    fabric_llpp0_araddr_s_o1	: out std_logic := '0';
    fabric_llpp0_araddr_s_o2	: out std_logic := '0';
    fabric_llpp0_araddr_s_o3	: out std_logic := '0';
    fabric_llpp0_araddr_s_o4	: out std_logic := '0';
    fabric_llpp0_araddr_s_o5	: out std_logic := '0';
    fabric_llpp0_araddr_s_o6	: out std_logic := '0';
    fabric_llpp0_araddr_s_o7	: out std_logic := '0';
    fabric_llpp0_araddr_s_o8	: out std_logic := '0';
    fabric_llpp0_araddr_s_o9	: out std_logic := '0';
    fabric_llpp0_araddr_s_o10	: out std_logic := '0';
    fabric_llpp0_araddr_s_o11	: out std_logic := '0';
    fabric_llpp0_araddr_s_o12	: out std_logic := '0';
    fabric_llpp0_araddr_s_o13	: out std_logic := '0';
    fabric_llpp0_araddr_s_o14	: out std_logic := '0';
    fabric_llpp0_araddr_s_o15	: out std_logic := '0';
    fabric_llpp0_araddr_s_o16	: out std_logic := '0';
    fabric_llpp0_araddr_s_o17	: out std_logic := '0';
    fabric_llpp0_araddr_s_o18	: out std_logic := '0';
    fabric_llpp0_araddr_s_o19	: out std_logic := '0';
    fabric_llpp0_araddr_s_o20	: out std_logic := '0';
    fabric_llpp0_araddr_s_o21	: out std_logic := '0';
    fabric_llpp0_araddr_s_o22	: out std_logic := '0';
    fabric_llpp0_araddr_s_o23	: out std_logic := '0';
    fabric_llpp0_araddr_s_o24	: out std_logic := '0';
    fabric_llpp0_araddr_s_o25	: out std_logic := '0';
    fabric_llpp0_araddr_s_o26	: out std_logic := '0';
    fabric_llpp0_araddr_s_o27	: out std_logic := '0';
    fabric_llpp0_araddr_s_o28	: out std_logic := '0';
    fabric_llpp0_araddr_s_o29	: out std_logic := '0';
    fabric_llpp0_araddr_s_o30	: out std_logic := '0';
    fabric_llpp0_araddr_s_o31	: out std_logic := '0';
    fabric_llpp0_araddr_s_o32	: out std_logic := '0';
    fabric_llpp0_arburst_s_o1	: out std_logic := '0';
    fabric_llpp0_arburst_s_o2	: out std_logic := '0';
    fabric_llpp0_arcache_s_o1	: out std_logic := '0';
    fabric_llpp0_arcache_s_o2	: out std_logic := '0';
    fabric_llpp0_arcache_s_o3	: out std_logic := '0';
    fabric_llpp0_arcache_s_o4	: out std_logic := '0';
    fabric_llpp0_arid_s_o1	: out std_logic := '0';
    fabric_llpp0_arid_s_o2	: out std_logic := '0';
    fabric_llpp0_arid_s_o3	: out std_logic := '0';
    fabric_llpp0_arid_s_o4	: out std_logic := '0';
    fabric_llpp0_arid_s_o5	: out std_logic := '0';
    fabric_llpp0_arid_s_o6	: out std_logic := '0';
    fabric_llpp0_arid_s_o7	: out std_logic := '0';
    fabric_llpp0_arid_s_o8	: out std_logic := '0';
    fabric_llpp0_arid_s_o9	: out std_logic := '0';
    fabric_llpp0_arid_s_o10	: out std_logic := '0';
    fabric_llpp0_arid_s_o11	: out std_logic := '0';
    fabric_llpp0_arid_s_o12	: out std_logic := '0';
    fabric_llpp0_arlen_s_o1	: out std_logic := '0';
    fabric_llpp0_arlen_s_o2	: out std_logic := '0';
    fabric_llpp0_arlen_s_o3	: out std_logic := '0';
    fabric_llpp0_arlen_s_o4	: out std_logic := '0';
    fabric_llpp0_arlen_s_o5	: out std_logic := '0';
    fabric_llpp0_arlen_s_o6	: out std_logic := '0';
    fabric_llpp0_arlen_s_o7	: out std_logic := '0';
    fabric_llpp0_arlen_s_o8	: out std_logic := '0';
    fabric_llpp0_arlock_s_o	: out std_logic := '0';
    fabric_llpp0_arprot_s_o1	: out std_logic := '0';
    fabric_llpp0_arprot_s_o2	: out std_logic := '0';
    fabric_llpp0_arprot_s_o3	: out std_logic := '0';
    fabric_llpp0_arqos_s_o1	: out std_logic := '0';
    fabric_llpp0_arqos_s_o2	: out std_logic := '0';
    fabric_llpp0_arqos_s_o3	: out std_logic := '0';
    fabric_llpp0_arqos_s_o4	: out std_logic := '0';
    fabric_llpp0_arsize_s_o1	: out std_logic := '0';
    fabric_llpp0_arsize_s_o2	: out std_logic := '0';
    fabric_llpp0_arsize_s_o3	: out std_logic := '0';
    fabric_llpp0_arvalid_s_o	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o1	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o2	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o3	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o4	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o5	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o6	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o7	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o8	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o9	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o10	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o11	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o12	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o13	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o14	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o15	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o16	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o17	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o18	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o19	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o20	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o21	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o22	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o23	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o24	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o25	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o26	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o27	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o28	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o29	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o30	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o31	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o32	: out std_logic := '0';
    fabric_llpp0_awburst_s_o1	: out std_logic := '0';
    fabric_llpp0_awburst_s_o2	: out std_logic := '0';
    fabric_llpp0_awcache_s_o1	: out std_logic := '0';
    fabric_llpp0_awcache_s_o2	: out std_logic := '0';
    fabric_llpp0_awcache_s_o3	: out std_logic := '0';
    fabric_llpp0_awcache_s_o4	: out std_logic := '0';
    fabric_llpp0_awid_s_o1	: out std_logic := '0';
    fabric_llpp0_awid_s_o2	: out std_logic := '0';
    fabric_llpp0_awid_s_o3	: out std_logic := '0';
    fabric_llpp0_awid_s_o4	: out std_logic := '0';
    fabric_llpp0_awid_s_o5	: out std_logic := '0';
    fabric_llpp0_awid_s_o6	: out std_logic := '0';
    fabric_llpp0_awid_s_o7	: out std_logic := '0';
    fabric_llpp0_awid_s_o8	: out std_logic := '0';
    fabric_llpp0_awid_s_o9	: out std_logic := '0';
    fabric_llpp0_awid_s_o10	: out std_logic := '0';
    fabric_llpp0_awid_s_o11	: out std_logic := '0';
    fabric_llpp0_awid_s_o12	: out std_logic := '0';
    fabric_llpp0_awlen_s_o1	: out std_logic := '0';
    fabric_llpp0_awlen_s_o2	: out std_logic := '0';
    fabric_llpp0_awlen_s_o3	: out std_logic := '0';
    fabric_llpp0_awlen_s_o4	: out std_logic := '0';
    fabric_llpp0_awlen_s_o5	: out std_logic := '0';
    fabric_llpp0_awlen_s_o6	: out std_logic := '0';
    fabric_llpp0_awlen_s_o7	: out std_logic := '0';
    fabric_llpp0_awlen_s_o8	: out std_logic := '0';
    fabric_llpp0_awlock_s_o	: out std_logic := '0';
    fabric_llpp0_awprot_s_o1	: out std_logic := '0';
    fabric_llpp0_awprot_s_o2	: out std_logic := '0';
    fabric_llpp0_awprot_s_o3	: out std_logic := '0';
    fabric_llpp0_awqos_s_o1	: out std_logic := '0';
    fabric_llpp0_awqos_s_o2	: out std_logic := '0';
    fabric_llpp0_awqos_s_o3	: out std_logic := '0';
    fabric_llpp0_awqos_s_o4	: out std_logic := '0';
    fabric_llpp0_awsize_s_o1	: out std_logic := '0';
    fabric_llpp0_awsize_s_o2	: out std_logic := '0';
    fabric_llpp0_awsize_s_o3	: out std_logic := '0';
    fabric_llpp0_awvalid_s_o	: out std_logic := '0';
    fabric_llpp0_bready_s_o	: out std_logic := '0';
    fabric_llpp0_rready_s_o	: out std_logic := '0';
    fabric_llpp0_wdata_s_o1	: out std_logic := '0';
    fabric_llpp0_wdata_s_o2	: out std_logic := '0';
    fabric_llpp0_wdata_s_o3	: out std_logic := '0';
    fabric_llpp0_wdata_s_o4	: out std_logic := '0';
    fabric_llpp0_wdata_s_o5	: out std_logic := '0';
    fabric_llpp0_wdata_s_o6	: out std_logic := '0';
    fabric_llpp0_wdata_s_o7	: out std_logic := '0';
    fabric_llpp0_wdata_s_o8	: out std_logic := '0';
    fabric_llpp0_wdata_s_o9	: out std_logic := '0';
    fabric_llpp0_wdata_s_o10	: out std_logic := '0';
    fabric_llpp0_wdata_s_o11	: out std_logic := '0';
    fabric_llpp0_wdata_s_o12	: out std_logic := '0';
    fabric_llpp0_wdata_s_o13	: out std_logic := '0';
    fabric_llpp0_wdata_s_o14	: out std_logic := '0';
    fabric_llpp0_wdata_s_o15	: out std_logic := '0';
    fabric_llpp0_wdata_s_o16	: out std_logic := '0';
    fabric_llpp0_wdata_s_o17	: out std_logic := '0';
    fabric_llpp0_wdata_s_o18	: out std_logic := '0';
    fabric_llpp0_wdata_s_o19	: out std_logic := '0';
    fabric_llpp0_wdata_s_o20	: out std_logic := '0';
    fabric_llpp0_wdata_s_o21	: out std_logic := '0';
    fabric_llpp0_wdata_s_o22	: out std_logic := '0';
    fabric_llpp0_wdata_s_o23	: out std_logic := '0';
    fabric_llpp0_wdata_s_o24	: out std_logic := '0';
    fabric_llpp0_wdata_s_o25	: out std_logic := '0';
    fabric_llpp0_wdata_s_o26	: out std_logic := '0';
    fabric_llpp0_wdata_s_o27	: out std_logic := '0';
    fabric_llpp0_wdata_s_o28	: out std_logic := '0';
    fabric_llpp0_wdata_s_o29	: out std_logic := '0';
    fabric_llpp0_wdata_s_o30	: out std_logic := '0';
    fabric_llpp0_wdata_s_o31	: out std_logic := '0';
    fabric_llpp0_wdata_s_o32	: out std_logic := '0';
    fabric_llpp0_wlast_s_o	: out std_logic := '0';
    fabric_llpp0_wstrb_s_o1	: out std_logic := '0';
    fabric_llpp0_wstrb_s_o2	: out std_logic := '0';
    fabric_llpp0_wstrb_s_o3	: out std_logic := '0';
    fabric_llpp0_wstrb_s_o4	: out std_logic := '0';
    fabric_llpp0_wvalid_s_o	: out std_logic := '0';
    fabric_llpp0_arready_s_i	: in std_logic := '0';
    fabric_llpp0_awready_s_i	: in std_logic := '0';
    fabric_llpp0_bid_s_i1	: in std_logic := '0';
    fabric_llpp0_bid_s_i2	: in std_logic := '0';
    fabric_llpp0_bid_s_i3	: in std_logic := '0';
    fabric_llpp0_bid_s_i4	: in std_logic := '0';
    fabric_llpp0_bid_s_i5	: in std_logic := '0';
    fabric_llpp0_bid_s_i6	: in std_logic := '0';
    fabric_llpp0_bid_s_i7	: in std_logic := '0';
    fabric_llpp0_bid_s_i8	: in std_logic := '0';
    fabric_llpp0_bid_s_i9	: in std_logic := '0';
    fabric_llpp0_bid_s_i10	: in std_logic := '0';
    fabric_llpp0_bid_s_i11	: in std_logic := '0';
    fabric_llpp0_bid_s_i12	: in std_logic := '0';
    fabric_llpp0_bresp_s_i1	: in std_logic := '0';
    fabric_llpp0_bresp_s_i2	: in std_logic := '0';
    fabric_llpp0_bvalid_s_i	: in std_logic := '0';
    fabric_llpp0_rdata_s_i1	: in std_logic := '0';
    fabric_llpp0_rdata_s_i2	: in std_logic := '0';
    fabric_llpp0_rdata_s_i3	: in std_logic := '0';
    fabric_llpp0_rdata_s_i4	: in std_logic := '0';
    fabric_llpp0_rdata_s_i5	: in std_logic := '0';
    fabric_llpp0_rdata_s_i6	: in std_logic := '0';
    fabric_llpp0_rdata_s_i7	: in std_logic := '0';
    fabric_llpp0_rdata_s_i8	: in std_logic := '0';
    fabric_llpp0_rdata_s_i9	: in std_logic := '0';
    fabric_llpp0_rdata_s_i10	: in std_logic := '0';
    fabric_llpp0_rdata_s_i11	: in std_logic := '0';
    fabric_llpp0_rdata_s_i12	: in std_logic := '0';
    fabric_llpp0_rdata_s_i13	: in std_logic := '0';
    fabric_llpp0_rdata_s_i14	: in std_logic := '0';
    fabric_llpp0_rdata_s_i15	: in std_logic := '0';
    fabric_llpp0_rdata_s_i16	: in std_logic := '0';
    fabric_llpp0_rdata_s_i17	: in std_logic := '0';
    fabric_llpp0_rdata_s_i18	: in std_logic := '0';
    fabric_llpp0_rdata_s_i19	: in std_logic := '0';
    fabric_llpp0_rdata_s_i20	: in std_logic := '0';
    fabric_llpp0_rdata_s_i21	: in std_logic := '0';
    fabric_llpp0_rdata_s_i22	: in std_logic := '0';
    fabric_llpp0_rdata_s_i23	: in std_logic := '0';
    fabric_llpp0_rdata_s_i24	: in std_logic := '0';
    fabric_llpp0_rdata_s_i25	: in std_logic := '0';
    fabric_llpp0_rdata_s_i26	: in std_logic := '0';
    fabric_llpp0_rdata_s_i27	: in std_logic := '0';
    fabric_llpp0_rdata_s_i28	: in std_logic := '0';
    fabric_llpp0_rdata_s_i29	: in std_logic := '0';
    fabric_llpp0_rdata_s_i30	: in std_logic := '0';
    fabric_llpp0_rdata_s_i31	: in std_logic := '0';
    fabric_llpp0_rdata_s_i32	: in std_logic := '0';
    fabric_llpp0_rid_s_i1	: in std_logic := '0';
    fabric_llpp0_rid_s_i2	: in std_logic := '0';
    fabric_llpp0_rid_s_i3	: in std_logic := '0';
    fabric_llpp0_rid_s_i4	: in std_logic := '0';
    fabric_llpp0_rid_s_i5	: in std_logic := '0';
    fabric_llpp0_rid_s_i6	: in std_logic := '0';
    fabric_llpp0_rid_s_i7	: in std_logic := '0';
    fabric_llpp0_rid_s_i8	: in std_logic := '0';
    fabric_llpp0_rid_s_i9	: in std_logic := '0';
    fabric_llpp0_rid_s_i10	: in std_logic := '0';
    fabric_llpp0_rid_s_i11	: in std_logic := '0';
    fabric_llpp0_rid_s_i12	: in std_logic := '0';
    fabric_llpp0_rlast_s_i	: in std_logic := '0';
    fabric_llpp0_rresp_s_i1	: in std_logic := '0';
    fabric_llpp0_rresp_s_i2	: in std_logic := '0';
    fabric_llpp0_rvalid_s_i	: in std_logic := '0';
    fabric_llpp0_wready_s_i	: in std_logic := '0';
    fabric_llpp1_araddr_s_o1	: out std_logic := '0';
    fabric_llpp1_araddr_s_o2	: out std_logic := '0';
    fabric_llpp1_araddr_s_o3	: out std_logic := '0';
    fabric_llpp1_araddr_s_o4	: out std_logic := '0';
    fabric_llpp1_araddr_s_o5	: out std_logic := '0';
    fabric_llpp1_araddr_s_o6	: out std_logic := '0';
    fabric_llpp1_araddr_s_o7	: out std_logic := '0';
    fabric_llpp1_araddr_s_o8	: out std_logic := '0';
    fabric_llpp1_araddr_s_o9	: out std_logic := '0';
    fabric_llpp1_araddr_s_o10	: out std_logic := '0';
    fabric_llpp1_araddr_s_o11	: out std_logic := '0';
    fabric_llpp1_araddr_s_o12	: out std_logic := '0';
    fabric_llpp1_araddr_s_o13	: out std_logic := '0';
    fabric_llpp1_araddr_s_o14	: out std_logic := '0';
    fabric_llpp1_araddr_s_o15	: out std_logic := '0';
    fabric_llpp1_araddr_s_o16	: out std_logic := '0';
    fabric_llpp1_araddr_s_o17	: out std_logic := '0';
    fabric_llpp1_araddr_s_o18	: out std_logic := '0';
    fabric_llpp1_araddr_s_o19	: out std_logic := '0';
    fabric_llpp1_araddr_s_o20	: out std_logic := '0';
    fabric_llpp1_araddr_s_o21	: out std_logic := '0';
    fabric_llpp1_araddr_s_o22	: out std_logic := '0';
    fabric_llpp1_araddr_s_o23	: out std_logic := '0';
    fabric_llpp1_araddr_s_o24	: out std_logic := '0';
    fabric_llpp1_araddr_s_o25	: out std_logic := '0';
    fabric_llpp1_araddr_s_o26	: out std_logic := '0';
    fabric_llpp1_araddr_s_o27	: out std_logic := '0';
    fabric_llpp1_araddr_s_o28	: out std_logic := '0';
    fabric_llpp1_araddr_s_o29	: out std_logic := '0';
    fabric_llpp1_araddr_s_o30	: out std_logic := '0';
    fabric_llpp1_araddr_s_o31	: out std_logic := '0';
    fabric_llpp1_araddr_s_o32	: out std_logic := '0';
    fabric_llpp1_arburst_s_o1	: out std_logic := '0';
    fabric_llpp1_arburst_s_o2	: out std_logic := '0';
    fabric_llpp1_arcache_s_o1	: out std_logic := '0';
    fabric_llpp1_arcache_s_o2	: out std_logic := '0';
    fabric_llpp1_arcache_s_o3	: out std_logic := '0';
    fabric_llpp1_arcache_s_o4	: out std_logic := '0';
    fabric_llpp1_arid_s_o1	: out std_logic := '0';
    fabric_llpp1_arid_s_o2	: out std_logic := '0';
    fabric_llpp1_arid_s_o3	: out std_logic := '0';
    fabric_llpp1_arid_s_o4	: out std_logic := '0';
    fabric_llpp1_arid_s_o5	: out std_logic := '0';
    fabric_llpp1_arid_s_o6	: out std_logic := '0';
    fabric_llpp1_arid_s_o7	: out std_logic := '0';
    fabric_llpp1_arid_s_o8	: out std_logic := '0';
    fabric_llpp1_arid_s_o9	: out std_logic := '0';
    fabric_llpp1_arid_s_o10	: out std_logic := '0';
    fabric_llpp1_arid_s_o11	: out std_logic := '0';
    fabric_llpp1_arid_s_o12	: out std_logic := '0';
    fabric_llpp1_arlen_s_o1	: out std_logic := '0';
    fabric_llpp1_arlen_s_o2	: out std_logic := '0';
    fabric_llpp1_arlen_s_o3	: out std_logic := '0';
    fabric_llpp1_arlen_s_o4	: out std_logic := '0';
    fabric_llpp1_arlen_s_o5	: out std_logic := '0';
    fabric_llpp1_arlen_s_o6	: out std_logic := '0';
    fabric_llpp1_arlen_s_o7	: out std_logic := '0';
    fabric_llpp1_arlen_s_o8	: out std_logic := '0';
    fabric_llpp1_arlock_s_o	: out std_logic := '0';
    fabric_llpp1_arprot_s_o1	: out std_logic := '0';
    fabric_llpp1_arprot_s_o2	: out std_logic := '0';
    fabric_llpp1_arprot_s_o3	: out std_logic := '0';
    fabric_llpp1_arqos_s1_o1	: out std_logic := '0';
    fabric_llpp1_arqos_s1_o2	: out std_logic := '0';
    fabric_llpp1_arqos_s1_o3	: out std_logic := '0';
    fabric_llpp1_arqos_s1_o4	: out std_logic := '0';
    fabric_llpp1_arsize_s_o1	: out std_logic := '0';
    fabric_llpp1_arsize_s_o2	: out std_logic := '0';
    fabric_llpp1_arsize_s_o3	: out std_logic := '0';
    fabric_llpp1_arvalid_s_o	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o1	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o2	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o3	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o4	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o5	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o6	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o7	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o8	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o9	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o10	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o11	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o12	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o13	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o14	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o15	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o16	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o17	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o18	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o19	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o20	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o21	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o22	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o23	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o24	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o25	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o26	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o27	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o28	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o29	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o30	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o31	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o32	: out std_logic := '0';
    fabric_llpp1_awburst_s_o1	: out std_logic := '0';
    fabric_llpp1_awburst_s_o2	: out std_logic := '0';
    fabric_llpp1_awcache_s_o1	: out std_logic := '0';
    fabric_llpp1_awcache_s_o2	: out std_logic := '0';
    fabric_llpp1_awcache_s_o3	: out std_logic := '0';
    fabric_llpp1_awcache_s_o4	: out std_logic := '0';
    fabric_llpp1_awid_s_o1	: out std_logic := '0';
    fabric_llpp1_awid_s_o2	: out std_logic := '0';
    fabric_llpp1_awid_s_o3	: out std_logic := '0';
    fabric_llpp1_awid_s_o4	: out std_logic := '0';
    fabric_llpp1_awid_s_o5	: out std_logic := '0';
    fabric_llpp1_awid_s_o6	: out std_logic := '0';
    fabric_llpp1_awid_s_o7	: out std_logic := '0';
    fabric_llpp1_awid_s_o8	: out std_logic := '0';
    fabric_llpp1_awid_s_o9	: out std_logic := '0';
    fabric_llpp1_awid_s_o10	: out std_logic := '0';
    fabric_llpp1_awid_s_o11	: out std_logic := '0';
    fabric_llpp1_awid_s_o12	: out std_logic := '0';
    fabric_llpp1_awlen_s_o1	: out std_logic := '0';
    fabric_llpp1_awlen_s_o2	: out std_logic := '0';
    fabric_llpp1_awlen_s_o3	: out std_logic := '0';
    fabric_llpp1_awlen_s_o4	: out std_logic := '0';
    fabric_llpp1_awlen_s_o5	: out std_logic := '0';
    fabric_llpp1_awlen_s_o6	: out std_logic := '0';
    fabric_llpp1_awlen_s_o7	: out std_logic := '0';
    fabric_llpp1_awlen_s_o8	: out std_logic := '0';
    fabric_llpp1_awlock_s_o	: out std_logic := '0';
    fabric_llpp1_awprot_s_o1	: out std_logic := '0';
    fabric_llpp1_awprot_s_o2	: out std_logic := '0';
    fabric_llpp1_awprot_s_o3	: out std_logic := '0';
    fabric_llpp1_awqos_s_o1	: out std_logic := '0';
    fabric_llpp1_awqos_s_o2	: out std_logic := '0';
    fabric_llpp1_awqos_s_o3	: out std_logic := '0';
    fabric_llpp1_awqos_s_o4	: out std_logic := '0';
    fabric_llpp1_awsize_s_o1	: out std_logic := '0';
    fabric_llpp1_awsize_s_o2	: out std_logic := '0';
    fabric_llpp1_awsize_s_o3	: out std_logic := '0';
    fabric_llpp1_awvalid_s_o	: out std_logic := '0';
    fabric_llpp1_bready_s_o	: out std_logic := '0';
    fabric_llpp1_rready_s_o	: out std_logic := '0';
    fabric_llpp1_wdata_s_o1	: out std_logic := '0';
    fabric_llpp1_wdata_s_o2	: out std_logic := '0';
    fabric_llpp1_wdata_s_o3	: out std_logic := '0';
    fabric_llpp1_wdata_s_o4	: out std_logic := '0';
    fabric_llpp1_wdata_s_o5	: out std_logic := '0';
    fabric_llpp1_wdata_s_o6	: out std_logic := '0';
    fabric_llpp1_wdata_s_o7	: out std_logic := '0';
    fabric_llpp1_wdata_s_o8	: out std_logic := '0';
    fabric_llpp1_wdata_s_o9	: out std_logic := '0';
    fabric_llpp1_wdata_s_o10	: out std_logic := '0';
    fabric_llpp1_wdata_s_o11	: out std_logic := '0';
    fabric_llpp1_wdata_s_o12	: out std_logic := '0';
    fabric_llpp1_wdata_s_o13	: out std_logic := '0';
    fabric_llpp1_wdata_s_o14	: out std_logic := '0';
    fabric_llpp1_wdata_s_o15	: out std_logic := '0';
    fabric_llpp1_wdata_s_o16	: out std_logic := '0';
    fabric_llpp1_wdata_s_o17	: out std_logic := '0';
    fabric_llpp1_wdata_s_o18	: out std_logic := '0';
    fabric_llpp1_wdata_s_o19	: out std_logic := '0';
    fabric_llpp1_wdata_s_o20	: out std_logic := '0';
    fabric_llpp1_wdata_s_o21	: out std_logic := '0';
    fabric_llpp1_wdata_s_o22	: out std_logic := '0';
    fabric_llpp1_wdata_s_o23	: out std_logic := '0';
    fabric_llpp1_wdata_s_o24	: out std_logic := '0';
    fabric_llpp1_wdata_s_o25	: out std_logic := '0';
    fabric_llpp1_wdata_s_o26	: out std_logic := '0';
    fabric_llpp1_wdata_s_o27	: out std_logic := '0';
    fabric_llpp1_wdata_s_o28	: out std_logic := '0';
    fabric_llpp1_wdata_s_o29	: out std_logic := '0';
    fabric_llpp1_wdata_s_o30	: out std_logic := '0';
    fabric_llpp1_wdata_s_o31	: out std_logic := '0';
    fabric_llpp1_wdata_s_o32	: out std_logic := '0';
    fabric_llpp1_wlast_s_o	: out std_logic := '0';
    fabric_llpp1_wstrb_s_o1	: out std_logic := '0';
    fabric_llpp1_wstrb_s_o2	: out std_logic := '0';
    fabric_llpp1_wstrb_s_o3	: out std_logic := '0';
    fabric_llpp1_wstrb_s_o4	: out std_logic := '0';
    fabric_llpp1_wvalid_s_o	: out std_logic := '0';
    fabric_llpp1_arready_s_i	: in std_logic := '0';
    fabric_llpp1_awready_s_i	: in std_logic := '0';
    fabric_llpp1_bid_s_i1	: in std_logic := '0';
    fabric_llpp1_bid_s_i2	: in std_logic := '0';
    fabric_llpp1_bid_s_i3	: in std_logic := '0';
    fabric_llpp1_bid_s_i4	: in std_logic := '0';
    fabric_llpp1_bid_s_i5	: in std_logic := '0';
    fabric_llpp1_bid_s_i6	: in std_logic := '0';
    fabric_llpp1_bid_s_i7	: in std_logic := '0';
    fabric_llpp1_bid_s_i8	: in std_logic := '0';
    fabric_llpp1_bid_s_i9	: in std_logic := '0';
    fabric_llpp1_bid_s_i10	: in std_logic := '0';
    fabric_llpp1_bid_s_i11	: in std_logic := '0';
    fabric_llpp1_bid_s_i12	: in std_logic := '0';
    fabric_llpp1_bresp_s_i1	: in std_logic := '0';
    fabric_llpp1_bresp_s_i2	: in std_logic := '0';
    fabric_llpp1_bvalid_s_i	: in std_logic := '0';
    fabric_llpp1_rdata_s_i1	: in std_logic := '0';
    fabric_llpp1_rdata_s_i2	: in std_logic := '0';
    fabric_llpp1_rdata_s_i3	: in std_logic := '0';
    fabric_llpp1_rdata_s_i4	: in std_logic := '0';
    fabric_llpp1_rdata_s_i5	: in std_logic := '0';
    fabric_llpp1_rdata_s_i6	: in std_logic := '0';
    fabric_llpp1_rdata_s_i7	: in std_logic := '0';
    fabric_llpp1_rdata_s_i8	: in std_logic := '0';
    fabric_llpp1_rdata_s_i9	: in std_logic := '0';
    fabric_llpp1_rdata_s_i10	: in std_logic := '0';
    fabric_llpp1_rdata_s_i11	: in std_logic := '0';
    fabric_llpp1_rdata_s_i12	: in std_logic := '0';
    fabric_llpp1_rdata_s_i13	: in std_logic := '0';
    fabric_llpp1_rdata_s_i14	: in std_logic := '0';
    fabric_llpp1_rdata_s_i15	: in std_logic := '0';
    fabric_llpp1_rdata_s_i16	: in std_logic := '0';
    fabric_llpp1_rdata_s_i17	: in std_logic := '0';
    fabric_llpp1_rdata_s_i18	: in std_logic := '0';
    fabric_llpp1_rdata_s_i19	: in std_logic := '0';
    fabric_llpp1_rdata_s_i20	: in std_logic := '0';
    fabric_llpp1_rdata_s_i21	: in std_logic := '0';
    fabric_llpp1_rdata_s_i22	: in std_logic := '0';
    fabric_llpp1_rdata_s_i23	: in std_logic := '0';
    fabric_llpp1_rdata_s_i24	: in std_logic := '0';
    fabric_llpp1_rdata_s_i25	: in std_logic := '0';
    fabric_llpp1_rdata_s_i26	: in std_logic := '0';
    fabric_llpp1_rdata_s_i27	: in std_logic := '0';
    fabric_llpp1_rdata_s_i28	: in std_logic := '0';
    fabric_llpp1_rdata_s_i29	: in std_logic := '0';
    fabric_llpp1_rdata_s_i30	: in std_logic := '0';
    fabric_llpp1_rdata_s_i31	: in std_logic := '0';
    fabric_llpp1_rdata_s_i32	: in std_logic := '0';
    fabric_llpp1_rid_s_i1	: in std_logic := '0';
    fabric_llpp1_rid_s_i2	: in std_logic := '0';
    fabric_llpp1_rid_s_i3	: in std_logic := '0';
    fabric_llpp1_rid_s_i4	: in std_logic := '0';
    fabric_llpp1_rid_s_i5	: in std_logic := '0';
    fabric_llpp1_rid_s_i6	: in std_logic := '0';
    fabric_llpp1_rid_s_i7	: in std_logic := '0';
    fabric_llpp1_rid_s_i8	: in std_logic := '0';
    fabric_llpp1_rid_s_i9	: in std_logic := '0';
    fabric_llpp1_rid_s_i10	: in std_logic := '0';
    fabric_llpp1_rid_s_i11	: in std_logic := '0';
    fabric_llpp1_rid_s_i12	: in std_logic := '0';
    fabric_llpp1_rlast_s_i	: in std_logic := '0';
    fabric_llpp1_rresp_s_i1	: in std_logic := '0';
    fabric_llpp1_rresp_s_i2	: in std_logic := '0';
    fabric_llpp1_rvalid_s_i	: in std_logic := '0';
    fabric_llpp1_wready_s_i	: in std_logic := '0';
    fabric_llpp2_araddr_s_o1	: out std_logic := '0';
    fabric_llpp2_araddr_s_o2	: out std_logic := '0';
    fabric_llpp2_araddr_s_o3	: out std_logic := '0';
    fabric_llpp2_araddr_s_o4	: out std_logic := '0';
    fabric_llpp2_araddr_s_o5	: out std_logic := '0';
    fabric_llpp2_araddr_s_o6	: out std_logic := '0';
    fabric_llpp2_araddr_s_o7	: out std_logic := '0';
    fabric_llpp2_araddr_s_o8	: out std_logic := '0';
    fabric_llpp2_araddr_s_o9	: out std_logic := '0';
    fabric_llpp2_araddr_s_o10	: out std_logic := '0';
    fabric_llpp2_araddr_s_o11	: out std_logic := '0';
    fabric_llpp2_araddr_s_o12	: out std_logic := '0';
    fabric_llpp2_araddr_s_o13	: out std_logic := '0';
    fabric_llpp2_araddr_s_o14	: out std_logic := '0';
    fabric_llpp2_araddr_s_o15	: out std_logic := '0';
    fabric_llpp2_araddr_s_o16	: out std_logic := '0';
    fabric_llpp2_araddr_s_o17	: out std_logic := '0';
    fabric_llpp2_araddr_s_o18	: out std_logic := '0';
    fabric_llpp2_araddr_s_o19	: out std_logic := '0';
    fabric_llpp2_araddr_s_o20	: out std_logic := '0';
    fabric_llpp2_araddr_s_o21	: out std_logic := '0';
    fabric_llpp2_araddr_s_o22	: out std_logic := '0';
    fabric_llpp2_araddr_s_o23	: out std_logic := '0';
    fabric_llpp2_araddr_s_o24	: out std_logic := '0';
    fabric_llpp2_araddr_s_o25	: out std_logic := '0';
    fabric_llpp2_araddr_s_o26	: out std_logic := '0';
    fabric_llpp2_araddr_s_o27	: out std_logic := '0';
    fabric_llpp2_araddr_s_o28	: out std_logic := '0';
    fabric_llpp2_araddr_s_o29	: out std_logic := '0';
    fabric_llpp2_araddr_s_o30	: out std_logic := '0';
    fabric_llpp2_araddr_s_o31	: out std_logic := '0';
    fabric_llpp2_araddr_s_o32	: out std_logic := '0';
    fabric_llpp2_arburst_s_o1	: out std_logic := '0';
    fabric_llpp2_arburst_s_o2	: out std_logic := '0';
    fabric_llpp2_arcache_s_o1	: out std_logic := '0';
    fabric_llpp2_arcache_s_o2	: out std_logic := '0';
    fabric_llpp2_arcache_s_o3	: out std_logic := '0';
    fabric_llpp2_arcache_s_o4	: out std_logic := '0';
    fabric_llpp2_arid_s_o1	: out std_logic := '0';
    fabric_llpp2_arid_s_o2	: out std_logic := '0';
    fabric_llpp2_arid_s_o3	: out std_logic := '0';
    fabric_llpp2_arid_s_o4	: out std_logic := '0';
    fabric_llpp2_arid_s_o5	: out std_logic := '0';
    fabric_llpp2_arid_s_o6	: out std_logic := '0';
    fabric_llpp2_arid_s_o7	: out std_logic := '0';
    fabric_llpp2_arid_s_o8	: out std_logic := '0';
    fabric_llpp2_arid_s_o9	: out std_logic := '0';
    fabric_llpp2_arid_s_o10	: out std_logic := '0';
    fabric_llpp2_arid_s_o11	: out std_logic := '0';
    fabric_llpp2_arid_s_o12	: out std_logic := '0';
    fabric_llpp2_arlen_s_o1	: out std_logic := '0';
    fabric_llpp2_arlen_s_o2	: out std_logic := '0';
    fabric_llpp2_arlen_s_o3	: out std_logic := '0';
    fabric_llpp2_arlen_s_o4	: out std_logic := '0';
    fabric_llpp2_arlen_s_o5	: out std_logic := '0';
    fabric_llpp2_arlen_s_o6	: out std_logic := '0';
    fabric_llpp2_arlen_s_o7	: out std_logic := '0';
    fabric_llpp2_arlen_s_o8	: out std_logic := '0';
    fabric_llpp2_arlock_s_o	: out std_logic := '0';
    fabric_llpp2_arprot_s_o1	: out std_logic := '0';
    fabric_llpp2_arprot_s_o2	: out std_logic := '0';
    fabric_llpp2_arprot_s_o3	: out std_logic := '0';
    fabric_llpp2_arqos_s_o1	: out std_logic := '0';
    fabric_llpp2_arqos_s_o2	: out std_logic := '0';
    fabric_llpp2_arqos_s_o3	: out std_logic := '0';
    fabric_llpp2_arqos_s_o4	: out std_logic := '0';
    fabric_llpp2_arsize_s_o1	: out std_logic := '0';
    fabric_llpp2_arsize_s_o2	: out std_logic := '0';
    fabric_llpp2_arsize_s_o3	: out std_logic := '0';
    fabric_llpp2_arvalid_s_o	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o1	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o2	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o3	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o4	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o5	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o6	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o7	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o8	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o9	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o10	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o11	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o12	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o13	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o14	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o15	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o16	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o17	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o18	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o19	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o20	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o21	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o22	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o23	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o24	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o25	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o26	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o27	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o28	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o29	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o30	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o31	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o32	: out std_logic := '0';
    fabric_llpp2_awburst_s_o1	: out std_logic := '0';
    fabric_llpp2_awburst_s_o2	: out std_logic := '0';
    fabric_llpp2_awcache_s_o1	: out std_logic := '0';
    fabric_llpp2_awcache_s_o2	: out std_logic := '0';
    fabric_llpp2_awcache_s_o3	: out std_logic := '0';
    fabric_llpp2_awcache_s_o4	: out std_logic := '0';
    fabric_llpp2_awid_s_o1	: out std_logic := '0';
    fabric_llpp2_awid_s_o2	: out std_logic := '0';
    fabric_llpp2_awid_s_o3	: out std_logic := '0';
    fabric_llpp2_awid_s_o4	: out std_logic := '0';
    fabric_llpp2_awid_s_o5	: out std_logic := '0';
    fabric_llpp2_awid_s_o6	: out std_logic := '0';
    fabric_llpp2_awid_s_o7	: out std_logic := '0';
    fabric_llpp2_awid_s_o8	: out std_logic := '0';
    fabric_llpp2_awid_s_o9	: out std_logic := '0';
    fabric_llpp2_awid_s_o10	: out std_logic := '0';
    fabric_llpp2_awid_s_o11	: out std_logic := '0';
    fabric_llpp2_awid_s_o12	: out std_logic := '0';
    fabric_llpp2_awlen_s_o1	: out std_logic := '0';
    fabric_llpp2_awlen_s_o2	: out std_logic := '0';
    fabric_llpp2_awlen_s_o3	: out std_logic := '0';
    fabric_llpp2_awlen_s_o4	: out std_logic := '0';
    fabric_llpp2_awlen_s_o5	: out std_logic := '0';
    fabric_llpp2_awlen_s_o6	: out std_logic := '0';
    fabric_llpp2_awlen_s_o7	: out std_logic := '0';
    fabric_llpp2_awlen_s_o8	: out std_logic := '0';
    fabric_llpp2_awlock_s_o	: out std_logic := '0';
    fabric_llpp2_awprot_s_o1	: out std_logic := '0';
    fabric_llpp2_awprot_s_o2	: out std_logic := '0';
    fabric_llpp2_awprot_s_o3	: out std_logic := '0';
    fabric_llpp2_awqos_s_o1	: out std_logic := '0';
    fabric_llpp2_awqos_s_o2	: out std_logic := '0';
    fabric_llpp2_awqos_s_o3	: out std_logic := '0';
    fabric_llpp2_awqos_s_o4	: out std_logic := '0';
    fabric_llpp2_awsize_s_o1	: out std_logic := '0';
    fabric_llpp2_awsize_s_o2	: out std_logic := '0';
    fabric_llpp2_awsize_s_o3	: out std_logic := '0';
    fabric_llpp2_awvalid_s_o	: out std_logic := '0';
    fabric_llpp2_bready_s_o	: out std_logic := '0';
    fabric_llpp2_rready_s_o	: out std_logic := '0';
    fabric_llpp2_wdata_s_o1	: out std_logic := '0';
    fabric_llpp2_wdata_s_o2	: out std_logic := '0';
    fabric_llpp2_wdata_s_o3	: out std_logic := '0';
    fabric_llpp2_wdata_s_o4	: out std_logic := '0';
    fabric_llpp2_wdata_s_o5	: out std_logic := '0';
    fabric_llpp2_wdata_s_o6	: out std_logic := '0';
    fabric_llpp2_wdata_s_o7	: out std_logic := '0';
    fabric_llpp2_wdata_s_o8	: out std_logic := '0';
    fabric_llpp2_wdata_s_o9	: out std_logic := '0';
    fabric_llpp2_wdata_s_o10	: out std_logic := '0';
    fabric_llpp2_wdata_s_o11	: out std_logic := '0';
    fabric_llpp2_wdata_s_o12	: out std_logic := '0';
    fabric_llpp2_wdata_s_o13	: out std_logic := '0';
    fabric_llpp2_wdata_s_o14	: out std_logic := '0';
    fabric_llpp2_wdata_s_o15	: out std_logic := '0';
    fabric_llpp2_wdata_s_o16	: out std_logic := '0';
    fabric_llpp2_wdata_s_o17	: out std_logic := '0';
    fabric_llpp2_wdata_s_o18	: out std_logic := '0';
    fabric_llpp2_wdata_s_o19	: out std_logic := '0';
    fabric_llpp2_wdata_s_o20	: out std_logic := '0';
    fabric_llpp2_wdata_s_o21	: out std_logic := '0';
    fabric_llpp2_wdata_s_o22	: out std_logic := '0';
    fabric_llpp2_wdata_s_o23	: out std_logic := '0';
    fabric_llpp2_wdata_s_o24	: out std_logic := '0';
    fabric_llpp2_wdata_s_o25	: out std_logic := '0';
    fabric_llpp2_wdata_s_o26	: out std_logic := '0';
    fabric_llpp2_wdata_s_o27	: out std_logic := '0';
    fabric_llpp2_wdata_s_o28	: out std_logic := '0';
    fabric_llpp2_wdata_s_o29	: out std_logic := '0';
    fabric_llpp2_wdata_s_o30	: out std_logic := '0';
    fabric_llpp2_wdata_s_o31	: out std_logic := '0';
    fabric_llpp2_wdata_s_o32	: out std_logic := '0';
    fabric_llpp2_wlast_s_o	: out std_logic := '0';
    fabric_llpp2_wstrb_s_o1	: out std_logic := '0';
    fabric_llpp2_wstrb_s_o2	: out std_logic := '0';
    fabric_llpp2_wstrb_s_o3	: out std_logic := '0';
    fabric_llpp2_wstrb_s_o4	: out std_logic := '0';
    fabric_llpp2_wvalid_s_o	: out std_logic := '0';
    fabric_llpp2_arready_s_i	: in std_logic := '0';
    fabric_llpp2_awready_s_i	: in std_logic := '0';
    fabric_llpp2_bid_s_i1	: in std_logic := '0';
    fabric_llpp2_bid_s_i2	: in std_logic := '0';
    fabric_llpp2_bid_s_i3	: in std_logic := '0';
    fabric_llpp2_bid_s_i4	: in std_logic := '0';
    fabric_llpp2_bid_s_i5	: in std_logic := '0';
    fabric_llpp2_bid_s_i6	: in std_logic := '0';
    fabric_llpp2_bid_s_i7	: in std_logic := '0';
    fabric_llpp2_bid_s_i8	: in std_logic := '0';
    fabric_llpp2_bid_s_i9	: in std_logic := '0';
    fabric_llpp2_bid_s_i10	: in std_logic := '0';
    fabric_llpp2_bid_s_i11	: in std_logic := '0';
    fabric_llpp2_bid_s_i12	: in std_logic := '0';
    fabric_llpp2_bresp_s_i1	: in std_logic := '0';
    fabric_llpp2_bresp_s_i2	: in std_logic := '0';
    fabric_llpp2_bvalid_s_i	: in std_logic := '0';
    fabric_llpp2_rdata_s_i1	: in std_logic := '0';
    fabric_llpp2_rdata_s_i2	: in std_logic := '0';
    fabric_llpp2_rdata_s_i3	: in std_logic := '0';
    fabric_llpp2_rdata_s_i4	: in std_logic := '0';
    fabric_llpp2_rdata_s_i5	: in std_logic := '0';
    fabric_llpp2_rdata_s_i6	: in std_logic := '0';
    fabric_llpp2_rdata_s_i7	: in std_logic := '0';
    fabric_llpp2_rdata_s_i8	: in std_logic := '0';
    fabric_llpp2_rdata_s_i9	: in std_logic := '0';
    fabric_llpp2_rdata_s_i10	: in std_logic := '0';
    fabric_llpp2_rdata_s_i11	: in std_logic := '0';
    fabric_llpp2_rdata_s_i12	: in std_logic := '0';
    fabric_llpp2_rdata_s_i13	: in std_logic := '0';
    fabric_llpp2_rdata_s_i14	: in std_logic := '0';
    fabric_llpp2_rdata_s_i15	: in std_logic := '0';
    fabric_llpp2_rdata_s_i16	: in std_logic := '0';
    fabric_llpp2_rdata_s_i17	: in std_logic := '0';
    fabric_llpp2_rdata_s_i18	: in std_logic := '0';
    fabric_llpp2_rdata_s_i19	: in std_logic := '0';
    fabric_llpp2_rdata_s_i20	: in std_logic := '0';
    fabric_llpp2_rdata_s_i21	: in std_logic := '0';
    fabric_llpp2_rdata_s_i22	: in std_logic := '0';
    fabric_llpp2_rdata_s_i23	: in std_logic := '0';
    fabric_llpp2_rdata_s_i24	: in std_logic := '0';
    fabric_llpp2_rdata_s_i25	: in std_logic := '0';
    fabric_llpp2_rdata_s_i26	: in std_logic := '0';
    fabric_llpp2_rdata_s_i27	: in std_logic := '0';
    fabric_llpp2_rdata_s_i28	: in std_logic := '0';
    fabric_llpp2_rdata_s_i29	: in std_logic := '0';
    fabric_llpp2_rdata_s_i30	: in std_logic := '0';
    fabric_llpp2_rdata_s_i31	: in std_logic := '0';
    fabric_llpp2_rdata_s_i32	: in std_logic := '0';
    fabric_llpp2_rid_s_i1	: in std_logic := '0';
    fabric_llpp2_rid_s_i2	: in std_logic := '0';
    fabric_llpp2_rid_s_i3	: in std_logic := '0';
    fabric_llpp2_rid_s_i4	: in std_logic := '0';
    fabric_llpp2_rid_s_i5	: in std_logic := '0';
    fabric_llpp2_rid_s_i6	: in std_logic := '0';
    fabric_llpp2_rid_s_i7	: in std_logic := '0';
    fabric_llpp2_rid_s_i8	: in std_logic := '0';
    fabric_llpp2_rid_s_i9	: in std_logic := '0';
    fabric_llpp2_rid_s_i10	: in std_logic := '0';
    fabric_llpp2_rid_s_i11	: in std_logic := '0';
    fabric_llpp2_rid_s_i12	: in std_logic := '0';
    fabric_llpp2_rlast_s_i	: in std_logic := '0';
    fabric_llpp2_rresp_s_i1	: in std_logic := '0';
    fabric_llpp2_rresp_s_i2	: in std_logic := '0';
    fabric_llpp2_rvalid_s_i	: in std_logic := '0';
    fabric_llpp2_wready_s_i	: in std_logic := '0';
    fabric_llpp3_araddr_s_o1	: out std_logic := '0';
    fabric_llpp3_araddr_s_o2	: out std_logic := '0';
    fabric_llpp3_araddr_s_o3	: out std_logic := '0';
    fabric_llpp3_araddr_s_o4	: out std_logic := '0';
    fabric_llpp3_araddr_s_o5	: out std_logic := '0';
    fabric_llpp3_araddr_s_o6	: out std_logic := '0';
    fabric_llpp3_araddr_s_o7	: out std_logic := '0';
    fabric_llpp3_araddr_s_o8	: out std_logic := '0';
    fabric_llpp3_araddr_s_o9	: out std_logic := '0';
    fabric_llpp3_araddr_s_o10	: out std_logic := '0';
    fabric_llpp3_araddr_s_o11	: out std_logic := '0';
    fabric_llpp3_araddr_s_o12	: out std_logic := '0';
    fabric_llpp3_araddr_s_o13	: out std_logic := '0';
    fabric_llpp3_araddr_s_o14	: out std_logic := '0';
    fabric_llpp3_araddr_s_o15	: out std_logic := '0';
    fabric_llpp3_araddr_s_o16	: out std_logic := '0';
    fabric_llpp3_araddr_s_o17	: out std_logic := '0';
    fabric_llpp3_araddr_s_o18	: out std_logic := '0';
    fabric_llpp3_araddr_s_o19	: out std_logic := '0';
    fabric_llpp3_araddr_s_o20	: out std_logic := '0';
    fabric_llpp3_araddr_s_o21	: out std_logic := '0';
    fabric_llpp3_araddr_s_o22	: out std_logic := '0';
    fabric_llpp3_araddr_s_o23	: out std_logic := '0';
    fabric_llpp3_araddr_s_o24	: out std_logic := '0';
    fabric_llpp3_araddr_s_o25	: out std_logic := '0';
    fabric_llpp3_araddr_s_o26	: out std_logic := '0';
    fabric_llpp3_araddr_s_o27	: out std_logic := '0';
    fabric_llpp3_araddr_s_o28	: out std_logic := '0';
    fabric_llpp3_araddr_s_o29	: out std_logic := '0';
    fabric_llpp3_araddr_s_o30	: out std_logic := '0';
    fabric_llpp3_araddr_s_o31	: out std_logic := '0';
    fabric_llpp3_araddr_s_o32	: out std_logic := '0';
    fabric_llpp3_arburst_s_o1	: out std_logic := '0';
    fabric_llpp3_arburst_s_o2	: out std_logic := '0';
    fabric_llpp3_arcache_s_o1	: out std_logic := '0';
    fabric_llpp3_arcache_s_o2	: out std_logic := '0';
    fabric_llpp3_arcache_s_o3	: out std_logic := '0';
    fabric_llpp3_arcache_s_o4	: out std_logic := '0';
    fabric_llpp3_arid_s_o1	: out std_logic := '0';
    fabric_llpp3_arid_s_o2	: out std_logic := '0';
    fabric_llpp3_arid_s_o3	: out std_logic := '0';
    fabric_llpp3_arid_s_o4	: out std_logic := '0';
    fabric_llpp3_arid_s_o5	: out std_logic := '0';
    fabric_llpp3_arid_s_o6	: out std_logic := '0';
    fabric_llpp3_arid_s_o7	: out std_logic := '0';
    fabric_llpp3_arid_s_o8	: out std_logic := '0';
    fabric_llpp3_arid_s_o9	: out std_logic := '0';
    fabric_llpp3_arid_s_o10	: out std_logic := '0';
    fabric_llpp3_arid_s_o11	: out std_logic := '0';
    fabric_llpp3_arid_s_o12	: out std_logic := '0';
    fabric_llpp3_arlen_s_o1	: out std_logic := '0';
    fabric_llpp3_arlen_s_o2	: out std_logic := '0';
    fabric_llpp3_arlen_s_o3	: out std_logic := '0';
    fabric_llpp3_arlen_s_o4	: out std_logic := '0';
    fabric_llpp3_arlen_s_o5	: out std_logic := '0';
    fabric_llpp3_arlen_s_o6	: out std_logic := '0';
    fabric_llpp3_arlen_s_o7	: out std_logic := '0';
    fabric_llpp3_arlen_s_o8	: out std_logic := '0';
    fabric_llpp3_arlock_s_o	: out std_logic := '0';
    fabric_llpp3_arprot_s_o1	: out std_logic := '0';
    fabric_llpp3_arprot_s_o2	: out std_logic := '0';
    fabric_llpp3_arprot_s_o3	: out std_logic := '0';
    fabric_llpp3_arqos_s_o1	: out std_logic := '0';
    fabric_llpp3_arqos_s_o2	: out std_logic := '0';
    fabric_llpp3_arqos_s_o3	: out std_logic := '0';
    fabric_llpp3_arqos_s_o4	: out std_logic := '0';
    fabric_llpp3_arsize_s_o1	: out std_logic := '0';
    fabric_llpp3_arsize_s_o2	: out std_logic := '0';
    fabric_llpp3_arsize_s_o3	: out std_logic := '0';
    fabric_llpp3_arvalid_s_o	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o1	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o2	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o3	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o4	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o5	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o6	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o7	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o8	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o9	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o10	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o11	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o12	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o13	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o14	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o15	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o16	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o17	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o18	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o19	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o20	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o21	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o22	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o23	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o24	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o25	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o26	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o27	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o28	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o29	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o30	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o31	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o32	: out std_logic := '0';
    fabric_llpp3_awburst_s_o1	: out std_logic := '0';
    fabric_llpp3_awburst_s_o2	: out std_logic := '0';
    fabric_llpp3_awcache_s_o1	: out std_logic := '0';
    fabric_llpp3_awcache_s_o2	: out std_logic := '0';
    fabric_llpp3_awcache_s_o3	: out std_logic := '0';
    fabric_llpp3_awcache_s_o4	: out std_logic := '0';
    fabric_llpp3_awid_s_o1	: out std_logic := '0';
    fabric_llpp3_awid_s_o2	: out std_logic := '0';
    fabric_llpp3_awid_s_o3	: out std_logic := '0';
    fabric_llpp3_awid_s_o4	: out std_logic := '0';
    fabric_llpp3_awid_s_o5	: out std_logic := '0';
    fabric_llpp3_awid_s_o6	: out std_logic := '0';
    fabric_llpp3_awid_s_o7	: out std_logic := '0';
    fabric_llpp3_awid_s_o8	: out std_logic := '0';
    fabric_llpp3_awid_s_o9	: out std_logic := '0';
    fabric_llpp3_awid_s_o10	: out std_logic := '0';
    fabric_llpp3_awid_s_o11	: out std_logic := '0';
    fabric_llpp3_awid_s_o12	: out std_logic := '0';
    fabric_llpp3_awlen_s_o1	: out std_logic := '0';
    fabric_llpp3_awlen_s_o2	: out std_logic := '0';
    fabric_llpp3_awlen_s_o3	: out std_logic := '0';
    fabric_llpp3_awlen_s_o4	: out std_logic := '0';
    fabric_llpp3_awlen_s_o5	: out std_logic := '0';
    fabric_llpp3_awlen_s_o6	: out std_logic := '0';
    fabric_llpp3_awlen_s_o7	: out std_logic := '0';
    fabric_llpp3_awlen_s_o8	: out std_logic := '0';
    fabric_llpp3_awlock_s_o	: out std_logic := '0';
    fabric_llpp3_awprot_s_o1	: out std_logic := '0';
    fabric_llpp3_awprot_s_o2	: out std_logic := '0';
    fabric_llpp3_awprot_s_o3	: out std_logic := '0';
    fabric_llpp3_awqos_s_o1	: out std_logic := '0';
    fabric_llpp3_awqos_s_o2	: out std_logic := '0';
    fabric_llpp3_awqos_s_o3	: out std_logic := '0';
    fabric_llpp3_awqos_s_o4	: out std_logic := '0';
    fabric_llpp3_awsize_s_o1	: out std_logic := '0';
    fabric_llpp3_awsize_s_o2	: out std_logic := '0';
    fabric_llpp3_awsize_s_o3	: out std_logic := '0';
    fabric_llpp3_awvalid_s_o	: out std_logic := '0';
    fabric_llpp3_bready_s_o	: out std_logic := '0';
    fabric_llpp3_rready_s_o	: out std_logic := '0';
    fabric_llpp3_wdata_s_o1	: out std_logic := '0';
    fabric_llpp3_wdata_s_o2	: out std_logic := '0';
    fabric_llpp3_wdata_s_o3	: out std_logic := '0';
    fabric_llpp3_wdata_s_o4	: out std_logic := '0';
    fabric_llpp3_wdata_s_o5	: out std_logic := '0';
    fabric_llpp3_wdata_s_o6	: out std_logic := '0';
    fabric_llpp3_wdata_s_o7	: out std_logic := '0';
    fabric_llpp3_wdata_s_o8	: out std_logic := '0';
    fabric_llpp3_wdata_s_o9	: out std_logic := '0';
    fabric_llpp3_wdata_s_o10	: out std_logic := '0';
    fabric_llpp3_wdata_s_o11	: out std_logic := '0';
    fabric_llpp3_wdata_s_o12	: out std_logic := '0';
    fabric_llpp3_wdata_s_o13	: out std_logic := '0';
    fabric_llpp3_wdata_s_o14	: out std_logic := '0';
    fabric_llpp3_wdata_s_o15	: out std_logic := '0';
    fabric_llpp3_wdata_s_o16	: out std_logic := '0';
    fabric_llpp3_wdata_s_o17	: out std_logic := '0';
    fabric_llpp3_wdata_s_o18	: out std_logic := '0';
    fabric_llpp3_wdata_s_o19	: out std_logic := '0';
    fabric_llpp3_wdata_s_o20	: out std_logic := '0';
    fabric_llpp3_wdata_s_o21	: out std_logic := '0';
    fabric_llpp3_wdata_s_o22	: out std_logic := '0';
    fabric_llpp3_wdata_s_o23	: out std_logic := '0';
    fabric_llpp3_wdata_s_o24	: out std_logic := '0';
    fabric_llpp3_wdata_s_o25	: out std_logic := '0';
    fabric_llpp3_wdata_s_o26	: out std_logic := '0';
    fabric_llpp3_wdata_s_o27	: out std_logic := '0';
    fabric_llpp3_wdata_s_o28	: out std_logic := '0';
    fabric_llpp3_wdata_s_o29	: out std_logic := '0';
    fabric_llpp3_wdata_s_o30	: out std_logic := '0';
    fabric_llpp3_wdata_s_o31	: out std_logic := '0';
    fabric_llpp3_wdata_s_o32	: out std_logic := '0';
    fabric_llpp3_wlast_s_o	: out std_logic := '0';
    fabric_llpp3_wstrb_s_o1	: out std_logic := '0';
    fabric_llpp3_wstrb_s_o2	: out std_logic := '0';
    fabric_llpp3_wstrb_s_o3	: out std_logic := '0';
    fabric_llpp3_wstrb_s_o4	: out std_logic := '0';
    fabric_llpp3_wvalid_s_o	: out std_logic := '0';
    fabric_llpp3_arready_s_i	: in std_logic := '0';
    fabric_llpp3_awready_s_i	: in std_logic := '0';
    fabric_llpp3_bid_s_i1	: in std_logic := '0';
    fabric_llpp3_bid_s_i2	: in std_logic := '0';
    fabric_llpp3_bid_s_i3	: in std_logic := '0';
    fabric_llpp3_bid_s_i4	: in std_logic := '0';
    fabric_llpp3_bid_s_i5	: in std_logic := '0';
    fabric_llpp3_bid_s_i6	: in std_logic := '0';
    fabric_llpp3_bid_s_i7	: in std_logic := '0';
    fabric_llpp3_bid_s_i8	: in std_logic := '0';
    fabric_llpp3_bid_s_i9	: in std_logic := '0';
    fabric_llpp3_bid_s_i10	: in std_logic := '0';
    fabric_llpp3_bid_s_i11	: in std_logic := '0';
    fabric_llpp3_bid_s_i12	: in std_logic := '0';
    fabric_llpp3_bresp_s_i1	: in std_logic := '0';
    fabric_llpp3_bresp_s_i2	: in std_logic := '0';
    fabric_llpp3_bvalid_s_i	: in std_logic := '0';
    fabric_llpp3_rdata_s_i1	: in std_logic := '0';
    fabric_llpp3_rdata_s_i2	: in std_logic := '0';
    fabric_llpp3_rdata_s_i3	: in std_logic := '0';
    fabric_llpp3_rdata_s_i4	: in std_logic := '0';
    fabric_llpp3_rdata_s_i5	: in std_logic := '0';
    fabric_llpp3_rdata_s_i6	: in std_logic := '0';
    fabric_llpp3_rdata_s_i7	: in std_logic := '0';
    fabric_llpp3_rdata_s_i8	: in std_logic := '0';
    fabric_llpp3_rdata_s_i9	: in std_logic := '0';
    fabric_llpp3_rdata_s_i10	: in std_logic := '0';
    fabric_llpp3_rdata_s_i11	: in std_logic := '0';
    fabric_llpp3_rdata_s_i12	: in std_logic := '0';
    fabric_llpp3_rdata_s_i13	: in std_logic := '0';
    fabric_llpp3_rdata_s_i14	: in std_logic := '0';
    fabric_llpp3_rdata_s_i15	: in std_logic := '0';
    fabric_llpp3_rdata_s_i16	: in std_logic := '0';
    fabric_llpp3_rdata_s_i17	: in std_logic := '0';
    fabric_llpp3_rdata_s_i18	: in std_logic := '0';
    fabric_llpp3_rdata_s_i19	: in std_logic := '0';
    fabric_llpp3_rdata_s_i20	: in std_logic := '0';
    fabric_llpp3_rdata_s_i21	: in std_logic := '0';
    fabric_llpp3_rdata_s_i22	: in std_logic := '0';
    fabric_llpp3_rdata_s_i23	: in std_logic := '0';
    fabric_llpp3_rdata_s_i24	: in std_logic := '0';
    fabric_llpp3_rdata_s_i25	: in std_logic := '0';
    fabric_llpp3_rdata_s_i26	: in std_logic := '0';
    fabric_llpp3_rdata_s_i27	: in std_logic := '0';
    fabric_llpp3_rdata_s_i28	: in std_logic := '0';
    fabric_llpp3_rdata_s_i29	: in std_logic := '0';
    fabric_llpp3_rdata_s_i30	: in std_logic := '0';
    fabric_llpp3_rdata_s_i31	: in std_logic := '0';
    fabric_llpp3_rdata_s_i32	: in std_logic := '0';
    fabric_llpp3_rid_s_i1	: in std_logic := '0';
    fabric_llpp3_rid_s_i2	: in std_logic := '0';
    fabric_llpp3_rid_s_i3	: in std_logic := '0';
    fabric_llpp3_rid_s_i4	: in std_logic := '0';
    fabric_llpp3_rid_s_i5	: in std_logic := '0';
    fabric_llpp3_rid_s_i6	: in std_logic := '0';
    fabric_llpp3_rid_s_i7	: in std_logic := '0';
    fabric_llpp3_rid_s_i8	: in std_logic := '0';
    fabric_llpp3_rid_s_i9	: in std_logic := '0';
    fabric_llpp3_rid_s_i10	: in std_logic := '0';
    fabric_llpp3_rid_s_i11	: in std_logic := '0';
    fabric_llpp3_rid_s_i12	: in std_logic := '0';
    fabric_llpp3_rlast_s_i	: in std_logic := '0';
    fabric_llpp3_rresp_s_i1	: in std_logic := '0';
    fabric_llpp3_rresp_s_i2	: in std_logic := '0';
    fabric_llpp3_rvalid_s_i	: in std_logic := '0';
    fabric_llpp3_wready_s_i	: in std_logic := '0';
    fabric_qos_pprdata_o1	: out std_logic := '0';
    fabric_qos_pprdata_o2	: out std_logic := '0';
    fabric_qos_pprdata_o3	: out std_logic := '0';
    fabric_qos_pprdata_o4	: out std_logic := '0';
    fabric_qos_pprdata_o5	: out std_logic := '0';
    fabric_qos_pprdata_o6	: out std_logic := '0';
    fabric_qos_pprdata_o7	: out std_logic := '0';
    fabric_qos_pprdata_o8	: out std_logic := '0';
    fabric_qos_pprdata_o9	: out std_logic := '0';
    fabric_qos_pprdata_o10	: out std_logic := '0';
    fabric_qos_pprdata_o11	: out std_logic := '0';
    fabric_qos_pprdata_o12	: out std_logic := '0';
    fabric_qos_pprdata_o13	: out std_logic := '0';
    fabric_qos_pprdata_o14	: out std_logic := '0';
    fabric_qos_pprdata_o15	: out std_logic := '0';
    fabric_qos_pprdata_o16	: out std_logic := '0';
    fabric_qos_pprdata_o17	: out std_logic := '0';
    fabric_qos_pprdata_o18	: out std_logic := '0';
    fabric_qos_pprdata_o19	: out std_logic := '0';
    fabric_qos_pprdata_o20	: out std_logic := '0';
    fabric_qos_pprdata_o21	: out std_logic := '0';
    fabric_qos_pprdata_o22	: out std_logic := '0';
    fabric_qos_pprdata_o23	: out std_logic := '0';
    fabric_qos_pprdata_o24	: out std_logic := '0';
    fabric_qos_pprdata_o25	: out std_logic := '0';
    fabric_qos_pprdata_o26	: out std_logic := '0';
    fabric_qos_pprdata_o27	: out std_logic := '0';
    fabric_qos_pprdata_o28	: out std_logic := '0';
    fabric_qos_pprdata_o29	: out std_logic := '0';
    fabric_qos_pprdata_o30	: out std_logic := '0';
    fabric_qos_pprdata_o31	: out std_logic := '0';
    fabric_qos_pprdata_o32	: out std_logic := '0';
    fabric_qos_ppready_o	: out std_logic := '0';
    fabric_qos_ppslverr_o	: out std_logic := '0';
    fabric_qos_pclk_i	: in std_logic := '0';
    fabric_qos_ppaddr_i1	: in std_logic := '0';
    fabric_qos_ppaddr_i2	: in std_logic := '0';
    fabric_qos_ppaddr_i3	: in std_logic := '0';
    fabric_qos_ppaddr_i4	: in std_logic := '0';
    fabric_qos_ppaddr_i5	: in std_logic := '0';
    fabric_qos_ppaddr_i6	: in std_logic := '0';
    fabric_qos_ppaddr_i7	: in std_logic := '0';
    fabric_qos_ppaddr_i8	: in std_logic := '0';
    fabric_qos_ppaddr_i9	: in std_logic := '0';
    fabric_qos_ppaddr_i10	: in std_logic := '0';
    fabric_qos_ppaddr_i11	: in std_logic := '0';
    fabric_qos_ppaddr_i12	: in std_logic := '0';
    fabric_qos_ppaddr_i13	: in std_logic := '0';
    fabric_qos_ppaddr_i14	: in std_logic := '0';
    fabric_qos_ppaddr_i15	: in std_logic := '0';
    fabric_qos_ppaddr_i16	: in std_logic := '0';
    fabric_qos_ppaddr_i17	: in std_logic := '0';
    fabric_qos_ppaddr_i18	: in std_logic := '0';
    fabric_qos_ppaddr_i19	: in std_logic := '0';
    fabric_qos_ppaddr_i20	: in std_logic := '0';
    fabric_qos_ppaddr_i21	: in std_logic := '0';
    fabric_qos_ppaddr_i22	: in std_logic := '0';
    fabric_qos_ppaddr_i23	: in std_logic := '0';
    fabric_qos_ppaddr_i24	: in std_logic := '0';
    fabric_qos_ppaddr_i25	: in std_logic := '0';
    fabric_qos_ppaddr_i26	: in std_logic := '0';
    fabric_qos_ppaddr_i27	: in std_logic := '0';
    fabric_qos_ppaddr_i28	: in std_logic := '0';
    fabric_qos_ppaddr_i29	: in std_logic := '0';
    fabric_qos_ppaddr_i30	: in std_logic := '0';
    fabric_qos_ppaddr_i31	: in std_logic := '0';
    fabric_qos_ppaddr_i32	: in std_logic := '0';
    fabric_qos_ppenable_i	: in std_logic := '0';
    fabric_qos_ppwdata_i1	: in std_logic := '0';
    fabric_qos_ppwdata_i2	: in std_logic := '0';
    fabric_qos_ppwdata_i3	: in std_logic := '0';
    fabric_qos_ppwdata_i4	: in std_logic := '0';
    fabric_qos_ppwdata_i5	: in std_logic := '0';
    fabric_qos_ppwdata_i6	: in std_logic := '0';
    fabric_qos_ppwdata_i7	: in std_logic := '0';
    fabric_qos_ppwdata_i8	: in std_logic := '0';
    fabric_qos_ppwdata_i9	: in std_logic := '0';
    fabric_qos_ppwdata_i10	: in std_logic := '0';
    fabric_qos_ppwdata_i11	: in std_logic := '0';
    fabric_qos_ppwdata_i12	: in std_logic := '0';
    fabric_qos_ppwdata_i13	: in std_logic := '0';
    fabric_qos_ppwdata_i14	: in std_logic := '0';
    fabric_qos_ppwdata_i15	: in std_logic := '0';
    fabric_qos_ppwdata_i16	: in std_logic := '0';
    fabric_qos_ppwdata_i17	: in std_logic := '0';
    fabric_qos_ppwdata_i18	: in std_logic := '0';
    fabric_qos_ppwdata_i19	: in std_logic := '0';
    fabric_qos_ppwdata_i20	: in std_logic := '0';
    fabric_qos_ppwdata_i21	: in std_logic := '0';
    fabric_qos_ppwdata_i22	: in std_logic := '0';
    fabric_qos_ppwdata_i23	: in std_logic := '0';
    fabric_qos_ppwdata_i24	: in std_logic := '0';
    fabric_qos_ppwdata_i25	: in std_logic := '0';
    fabric_qos_ppwdata_i26	: in std_logic := '0';
    fabric_qos_ppwdata_i27	: in std_logic := '0';
    fabric_qos_ppwdata_i28	: in std_logic := '0';
    fabric_qos_ppwdata_i29	: in std_logic := '0';
    fabric_qos_ppwdata_i30	: in std_logic := '0';
    fabric_qos_ppwdata_i31	: in std_logic := '0';
    fabric_qos_ppwdata_i32	: in std_logic := '0';
    fabric_qos_ppwrite_i	: in std_logic := '0';
    fabric_qos_presetn_i	: in std_logic := '0';
    fabric_qos_psel_i	: in std_logic := '0';
    fabric_tnd_hssl_flushin_o	: out std_logic := '0';
    fabric_tnd_hssl_trigin_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o1	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o2	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o3	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o4	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o5	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o6	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o7	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o8	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o9	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o10	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o11	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o12	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o13	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o14	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o15	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o16	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o17	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o18	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o19	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o20	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o21	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o22	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o23	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o24	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o25	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o26	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o27	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o28	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o29	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o30	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o31	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o32	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_penable_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_psel_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o1	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o2	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o3	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o4	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o5	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o6	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o7	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o8	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o9	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o10	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o11	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o12	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o13	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o14	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o15	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o16	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o17	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o18	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o19	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o20	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o21	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o22	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o23	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o24	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o25	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o26	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o27	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o28	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o29	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o30	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o31	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o32	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwrite_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_afvalid_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_atready_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_syncreq_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o1	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o2	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o3	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o4	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o5	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o6	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o7	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o8	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o9	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o10	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o11	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o12	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o13	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o14	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o15	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o16	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o17	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o18	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o19	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o20	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o21	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o22	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o23	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o24	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o25	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o26	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o27	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o28	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o29	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o30	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o31	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o32	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_penable_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_psel_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o1	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o2	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o3	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o4	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o5	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o6	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o7	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o8	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o9	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o10	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o11	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o12	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o13	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o14	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o15	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o16	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o17	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o18	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o19	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o20	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o21	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o22	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o23	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o24	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o25	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o26	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o27	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o28	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o29	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o30	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o31	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o32	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwrite_o	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_afready_o	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atbytes_o1	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atbytes_o2	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atbytes_o3	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atbytes_o4	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o1	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o2	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o3	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o4	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o5	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o6	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o7	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o8	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o9	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o10	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o11	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o12	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o13	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o14	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o15	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o16	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o17	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o18	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o19	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o20	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o21	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o22	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o23	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o24	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o25	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o26	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o27	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o28	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o29	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o30	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o31	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o32	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o33	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o34	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o35	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o36	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o37	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o38	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o39	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o40	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o41	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o42	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o43	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o44	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o45	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o46	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o47	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o48	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o49	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o50	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o51	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o52	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o53	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o54	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o55	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o56	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o57	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o58	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o59	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o60	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o61	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o62	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o63	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o64	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o65	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o66	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o67	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o68	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o69	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o70	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o71	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o72	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o73	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o74	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o75	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o76	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o77	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o78	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o79	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o80	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o81	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o82	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o83	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o84	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o85	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o86	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o87	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o88	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o89	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o90	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o91	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o92	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o93	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o94	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o95	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o96	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o97	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o98	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o99	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o100	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o101	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o102	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o103	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o104	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o105	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o106	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o107	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o108	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o109	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o110	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o111	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o112	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o113	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o114	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o115	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o116	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o117	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o118	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o119	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o120	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o121	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o122	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o123	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o124	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o125	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o126	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o127	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atdata_o128	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o1	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o2	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o3	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o4	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o5	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o6	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atid_o7	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atvalid_o	: out std_logic := '0';
    fabric_tnd_trace_clk_traceoutportintf_o	: out std_logic := '0';
    fabric_tnd_trace_ctl_traceoutportintf_o	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o1	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o2	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o3	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o4	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o5	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o6	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o7	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o8	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o9	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o10	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o11	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o12	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o13	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o14	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o15	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o16	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o17	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o18	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o19	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o20	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o21	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o22	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o23	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o24	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o25	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o26	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o27	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o28	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o29	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o30	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o31	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o32	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o1	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o2	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o3	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o4	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o5	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o6	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o7	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o8	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o9	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o10	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o11	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o12	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o13	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o14	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o15	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o16	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o17	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o18	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o19	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o20	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o21	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o22	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o23	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o24	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o25	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o26	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o27	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o28	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o29	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o30	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o31	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o32	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o33	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o34	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o35	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o36	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o37	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o38	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o39	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o40	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o41	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o42	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o43	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o44	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o45	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o46	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o47	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o48	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o49	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o50	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o51	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o52	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o53	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o54	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o55	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o56	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o57	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o58	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o59	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o60	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o61	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o62	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o63	: out std_logic := '0';
    fabric_tsvalue_tsgen_fpga_o64	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i1	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i2	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i3	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i4	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i5	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i6	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i7	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i8	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i9	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i10	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i11	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i12	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i13	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i14	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i15	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i16	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i17	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i18	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i19	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i20	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i21	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i22	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i23	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i24	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i25	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i26	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i27	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i28	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i29	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i30	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i31	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_prdata_i32	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_pready_i	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_pslverr_i	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_afready_i	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atbytes_i1	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atbytes_i2	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atbytes_i3	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atbytes_i4	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i1	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i2	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i3	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i4	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i5	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i6	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i7	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i8	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i9	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i10	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i11	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i12	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i13	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i14	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i15	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i16	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i17	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i18	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i19	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i20	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i21	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i22	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i23	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i24	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i25	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i26	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i27	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i28	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i29	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i30	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i31	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i32	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i33	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i34	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i35	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i36	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i37	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i38	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i39	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i40	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i41	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i42	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i43	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i44	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i45	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i46	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i47	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i48	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i49	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i50	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i51	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i52	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i53	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i54	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i55	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i56	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i57	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i58	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i59	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i60	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i61	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i62	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i63	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i64	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i65	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i66	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i67	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i68	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i69	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i70	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i71	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i72	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i73	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i74	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i75	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i76	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i77	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i78	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i79	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i80	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i81	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i82	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i83	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i84	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i85	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i86	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i87	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i88	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i89	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i90	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i91	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i92	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i93	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i94	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i95	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i96	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i97	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i98	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i99	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i100	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i101	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i102	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i103	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i104	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i105	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i106	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i107	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i108	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i109	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i110	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i111	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i112	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i113	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i114	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i115	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i116	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i117	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i118	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i119	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i120	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i121	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i122	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i123	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i124	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i125	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i126	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i127	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atdata_i128	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i1	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i2	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i3	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i4	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i5	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i6	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atid_i7	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atvalid_i	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i1	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i2	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i3	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i4	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i5	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i6	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i7	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i8	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i9	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i10	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i11	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i12	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i13	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i14	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i15	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i16	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i17	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i18	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i19	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i20	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i21	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i22	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i23	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i24	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i25	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i26	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i27	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i28	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i29	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i30	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i31	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i32	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_pready_i	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_pslverr_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_afvalid_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_atready_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_syncreq_i	: in std_logic := '0';
    fabric_watchdog0_signal_0_o	: out std_logic := '0';
    fabric_watchdog0_signal_1_o	: out std_logic := '0';
    fabric_watchdog1_signal_0_o	: out std_logic := '0';
    fabric_watchdog1_signal_1_o	: out std_logic := '0';
    fabric_watchdog2_signal_0_o	: out std_logic := '0';
    fabric_watchdog2_signal_1_o	: out std_logic := '0';
    fabric_watchdog3_signal_0_o	: out std_logic := '0';
    fabric_watchdog3_signal_1_o	: out std_logic := '0';
    fabric_tst_pll_lock_o1	: out std_logic := '0';
    fabric_tst_pll_lock_o2	: out std_logic := '0';
    fabric_tst_pll_lock_o3	: out std_logic := '0';
    fabric_tst_pll_lock_o4	: out std_logic := '0';
    fabric_tst_pll_lock_o5	: out std_logic := '0';
    fabric_tst_pll_lock_o6	: out std_logic := '0';
    fabric_tst_pll_lock_o7	: out std_logic := '0';
    fabric_soc_mon_sensor_alarm_o	: out std_logic := '0';
    fabric_erom_fpga_cpu0_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cs_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cs_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cs_deviceen_i	: in std_logic := '0';
    fabric_erom_fpga_cs_rst_n_i	: in std_logic := '0';
    fabric_erom_fpga_debug_en_i	: in std_logic := '0';
    fabric_enable_TMR_i1	: in std_logic := '1';
    fabric_enable_TMR_i2	: in std_logic := '1';
    fabric_enable_TMR_i3	: in std_logic := '1'
);
end component NX_SOC_INTERFACE;

component NX_SOC_INTERFACE_WRAP is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    -- dahlia <-> fabric
    fabric_lowskew_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_lowskew_i	: in std_logic_vector(9   downto 0) := (others => '0');
    fabric_fpga_nic_rstn_i	: in std_logic_vector(9   downto 0) := (others => '0');
    fabric_fpga_pmrstn_i	: in std_logic := '0';
    fabric_fpga_sysrstn_i	: in std_logic := '0';
    fabric_fpga_trigger_in_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_trigger_out_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_interrupt_in_i	: in std_logic_vector(119 downto 0) := (others => '0');
    fabric_sysc_hold_on_debug_i	: in std_logic := '0';
    fabric_fpga_events60_i	: in std_logic_vector(59  downto 0) := (others => '0');
    fabric_fpga_araddr_axi_s1_o	: out std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_arburst_axi_s1_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_arcache_axi_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arid_axi_s1_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_arlen_axi_s1_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_arlock_axi_s1_o	: out std_logic := '0';
    fabric_fpga_arprot_axi_s1_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arqos_axi_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arregion_axi_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arsize_axi_s1_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s1_o	: out std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_awburst_axi_s1_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_awcache_axi_s1_o	: out std_logic_vector(3  downto 0) := (others => '0');
    fabric_fpga_awid_axi_s1_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_awlen_axi_s1_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_awlock_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awprot_axi_s1_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awqos_axi_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awregion_axi_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awsize_axi_s1_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_bready_axi_s1_o	: out std_logic := '0';
    fabric_fpga_rready_axi_s1_o	: out std_logic := '0';
    fabric_fpga_wdata_axi_s1_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_wlast_axi_s1_o	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s1_o	: out std_logic_vector(15  downto 0) := (others => '0');
    fabric_fpga_wvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_awvalid_axi_s1_o	: out std_logic := '0';
    fabric_fpga_arready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_awready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_bid_axi_s1_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_bresp_axi_s1_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_bvalid_axi_s1_i	: in std_logic := '0';
    fabric_fpga_rdata_axi_s1_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_rid_axi_s1_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_rlast_axi_s1_i	: in std_logic := '0';
    fabric_fpga_rresp_axi_s1_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_rvalid_axi_s1_i	: in std_logic := '0';
    fabric_fpga_wready_axi_s1_i	: in std_logic := '0';
    fabric_fpga_araddr_axi_s2_o	: out std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_arburst_axi_s2_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_arcache_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arid_axi_s2_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_arlen_axi_s2_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_arlock_axi_s2_o	: out std_logic := '0';
    fabric_fpga_arprot_axi_s2_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arqos_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arregion_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arsize_axi_s2_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awaddr_axi_s2_o	: out std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_awburst_axi_s2_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_awcache_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awid_axi_s2_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_awlen_axi_s2_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_awlock_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awprot_axi_s2_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awqos_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awregion_axi_s2_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awsize_axi_s2_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_bready_axi_s2_o	: out std_logic := '0';
    fabric_fpga_rready_axi_s2_o	: out std_logic := '0';
    fabric_fpga_wdata_axi_s2_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_wlast_axi_s2_o	: out std_logic := '0';
    fabric_fpga_wstrb_axi_s2_o	: out std_logic_vector(15  downto 0) := (others => '0');
    fabric_fpga_wvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_awvalid_axi_s2_o	: out std_logic := '0';
    fabric_fpga_arready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_awready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_bid_axi_s2_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_bresp_axi_s2_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_bvalid_axi_s2_i	: in std_logic := '0';
    fabric_fpga_rdata_axi_s2_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_rid_axi_s2_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_fpga_rlast_axi_s2_i	: in std_logic := '0';
    fabric_fpga_rresp_axi_s2_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_rvalid_axi_s2_i	: in std_logic := '0';
    fabric_fpga_wready_axi_s2_i	: in std_logic := '0';
    fabric_fpga_arready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_awready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_bid_axi_m1_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_bresp_axi_m1_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_bvalid_axi_m1_o	: out std_logic := '0';
    fabric_fpga_dma_ack_m1_o	: out std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_finish_m1_o	: out std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_rdata_axi_m1_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_rid_axi_m1_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_rlast_axi_m1_o	: out std_logic := '0';
    fabric_fpga_rresp_axi_m1_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_rvalid_axi_m1_o	: out std_logic := '0';
    fabric_fpga_wready_axi_m1_o	: out std_logic := '0';
    fabric_fpga_araddr_axi_m1_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_arburst_axi_m1_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_arcache_axi_m1_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arid_axi_m1_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_arlen_axi_m1_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_arlock_axi_m1_i	: in std_logic := '0';
    fabric_fpga_arprot_axi_m1_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arqos_axi_m1_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arsize_axi_m1_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m1_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_awburst_axi_m1_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_awcache_axi_m1_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awid_axi_m1_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_awlen_axi_m1_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_awlock_axi_m1_i	: in std_logic := '0';
    fabric_fpga_awprot_axi_m1_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awqos_axi_m1_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awsize_axi_m1_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_bready_axi_m1_i	: in std_logic := '0';
    fabric_fpga_dma_last_m1_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_req_m1_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_single_m1_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_rready_axi_m1_i	: in std_logic := '0';
    fabric_fpga_wdata_axi_m1_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_wlast_axi_m1_i	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m1_i	: in std_logic_vector(15  downto 0) := (others => '0');
    fabric_fpga_wvalid_axi_m1_i	: in std_logic := '0';
    fabric_fpga_arready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_awready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_bid_axi_m2_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_bresp_axi_m2_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_bvalid_axi_m2_o	: out std_logic := '0';
    fabric_fpga_dma_ack_m2_o	: out std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_finish_m2_o	: out std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_rdata_axi_m2_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_rid_axi_m2_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_rlast_axi_m2_o	: out std_logic := '0';
    fabric_fpga_rresp_axi_m2_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_rvalid_axi_m2_o	: out std_logic := '0';
    fabric_fpga_wready_axi_m2_o	: out std_logic := '0';
    fabric_fpga_araddr_axi_m2_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_arburst_axi_m2_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_arcache_axi_m2_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arid_axi_m2_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_arlen_axi_m2_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_arlock_axi_m2_i	: in std_logic := '0';
    fabric_fpga_arprot_axi_m2_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arqos_axi_m2_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_arsize_axi_m2_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_arvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_awaddr_axi_m2_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_awburst_axi_m2_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_awcache_axi_m2_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awid_axi_m2_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_awlen_axi_m2_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_awlock_axi_m2_i	: in std_logic := '0';
    fabric_fpga_awprot_axi_m2_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awqos_axi_m2_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_awsize_axi_m2_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_awvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_bready_axi_m2_i	: in std_logic := '0';
    fabric_fpga_dma_last_m2_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_req_m2_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_dma_single_m2_i	: in std_logic_vector(5   downto 0) := (others => '0');
    fabric_fpga_rready_axi_m2_i	: in std_logic := '0';
    fabric_fpga_wdata_axi_m2_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_wlast_axi_m2_i	: in std_logic := '0';
    fabric_fpga_wstrb_axi_m2_i	: in std_logic_vector(15  downto 0) := (others => '0');
    fabric_fpga_wvalid_axi_m2_i	: in std_logic := '0';
    fabric_fpga_ddr0_arready_o	: out std_logic := '0';
    fabric_fpga_ddr0_awready_o	: out std_logic := '0';
    fabric_fpga_ddr0_bid_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_ddr0_bresp_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_ddr0_bvalid_o	: out std_logic := '0';
    fabric_fpga_ddr0_rdata_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_ddr0_rid_o	: out std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_ddr0_rlast_o	: out std_logic := '0';
    fabric_fpga_ddr0_rresp_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_ddr0_rvalid_o	: out std_logic := '0';
    fabric_fpga_ddr0_wready_o	: out std_logic := '0';
    fabric_fpga_ddr0_araddr_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_ddr0_arburst_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_ddr0_arcache_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_ddr0_arid_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_ddr0_arlen_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_ddr0_arlock_i	: in std_logic := '0';
    fabric_fpga_ddr0_arprot_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_ddr0_arqos_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_ddr0_arsize_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_ddr0_arvalid_i	: in std_logic := '0';
    fabric_fpga_ddr0_awaddr_i	: in std_logic_vector(39  downto 0) := (others => '0');
    fabric_fpga_ddr0_awburst_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_fpga_ddr0_awcache_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_ddr0_awid_i	: in std_logic_vector(4   downto 0) := (others => '0');
    fabric_fpga_ddr0_awlen_i	: in std_logic_vector(7   downto 0) := (others => '0');
    fabric_fpga_ddr0_awlock_i	: in std_logic := '0';
    fabric_fpga_ddr0_awprot_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_ddr0_awqos_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_fpga_ddr0_awsize_i	: in std_logic_vector(2   downto 0) := (others => '0');
    fabric_fpga_ddr0_awvalid_i	: in std_logic := '0';
    fabric_fpga_ddr0_bready_i	: in std_logic := '0';
    fabric_fpga_ddr0_rready_i	: in std_logic := '0';
    fabric_fpga_ddr0_wdata_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_fpga_ddr0_wlast_i	: in std_logic := '0';
    fabric_fpga_ddr0_wstrb_i	: in std_logic_vector(15  downto 0) := (others => '0');
    fabric_fpga_ddr0_wvalid_i	: in std_logic := '0';
    fabric_fpga_paddr_apb_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_fpga_penable_apb_o	: out std_logic := '0';
    fabric_fpga_psel_apb_o	: out std_logic := '0';
    fabric_fpga_pwdata_apb_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_fpga_pwrite_apb_o	: out std_logic := '0';
    fabric_fpga_prdata_apb_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_fpga_pready_apb_i	: in std_logic := '0';
    fabric_fpga_pslverr_apb_i	: in std_logic := '0';
    fabric_llpp0_araddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp0_arburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp0_arcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp0_arid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp0_arlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp0_arlock_s_o	: out std_logic := '0';
    fabric_llpp0_arprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp0_arqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp0_arsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp0_arvalid_s_o	: out std_logic := '0';
    fabric_llpp0_awaddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp0_awburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp0_awcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp0_awid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp0_awlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp0_awlock_s_o	: out std_logic := '0';
    fabric_llpp0_awprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp0_awqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp0_awsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp0_awvalid_s_o	: out std_logic := '0';
    fabric_llpp0_bready_s_o	: out std_logic := '0';
    fabric_llpp0_rready_s_o	: out std_logic := '0';
    fabric_llpp0_wdata_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp0_wlast_s_o	: out std_logic := '0';
    fabric_llpp0_wstrb_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp0_wvalid_s_o	: out std_logic := '0';
    fabric_llpp0_arready_s_i	: in std_logic := '0';
    fabric_llpp0_awready_s_i	: in std_logic := '0';
    fabric_llpp0_bid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp0_bresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp0_bvalid_s_i	: in std_logic := '0';
    fabric_llpp0_rdata_s_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp0_rid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp0_rlast_s_i	: in std_logic := '0';
    fabric_llpp0_rresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp0_rvalid_s_i	: in std_logic := '0';
    fabric_llpp0_wready_s_i	: in std_logic := '0';
    fabric_llpp1_araddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp1_arburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp1_arcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp1_arid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp1_arlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp1_arlock_s_o	: out std_logic := '0';
    fabric_llpp1_arprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp1_arqos_s1_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp1_arsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp1_arvalid_s_o	: out std_logic := '0';
    fabric_llpp1_awaddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp1_awburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp1_awcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp1_awid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp1_awlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp1_awlock_s_o	: out std_logic := '0';
    fabric_llpp1_awprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp1_awqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp1_awsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp1_awvalid_s_o	: out std_logic := '0';
    fabric_llpp1_bready_s_o	: out std_logic := '0';
    fabric_llpp1_rready_s_o	: out std_logic := '0';
    fabric_llpp1_wdata_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp1_wlast_s_o	: out std_logic := '0';
    fabric_llpp1_wstrb_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp1_wvalid_s_o	: out std_logic := '0';
    fabric_llpp1_arready_s_i	: in std_logic := '0';
    fabric_llpp1_awready_s_i	: in std_logic := '0';
    fabric_llpp1_bid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp1_bresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp1_bvalid_s_i	: in std_logic := '0';
    fabric_llpp1_rdata_s_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp1_rid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp1_rlast_s_i	: in std_logic := '0';
    fabric_llpp1_rresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp1_rvalid_s_i	: in std_logic := '0';
    fabric_llpp1_wready_s_i	: in std_logic := '0';
    fabric_llpp2_araddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp2_arburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp2_arcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp2_arid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp2_arlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp2_arlock_s_o	: out std_logic := '0';
    fabric_llpp2_arprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp2_arqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp2_arsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp2_arvalid_s_o	: out std_logic := '0';
    fabric_llpp2_awaddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp2_awburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp2_awcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp2_awid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp2_awlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp2_awlock_s_o	: out std_logic := '0';
    fabric_llpp2_awprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp2_awqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp2_awsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp2_awvalid_s_o	: out std_logic := '0';
    fabric_llpp2_bready_s_o	: out std_logic := '0';
    fabric_llpp2_rready_s_o	: out std_logic := '0';
    fabric_llpp2_wdata_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp2_wlast_s_o	: out std_logic := '0';
    fabric_llpp2_wstrb_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp2_wvalid_s_o	: out std_logic := '0';
    fabric_llpp2_arready_s_i	: in std_logic := '0';
    fabric_llpp2_awready_s_i	: in std_logic := '0';
    fabric_llpp2_bid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp2_bresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp2_bvalid_s_i	: in std_logic := '0';
    fabric_llpp2_rdata_s_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp2_rid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp2_rlast_s_i	: in std_logic := '0';
    fabric_llpp2_rresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp2_rvalid_s_i	: in std_logic := '0';
    fabric_llpp2_wready_s_i	: in std_logic := '0';
    fabric_llpp3_araddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp3_arburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp3_arcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp3_arid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp3_arlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp3_arlock_s_o	: out std_logic := '0';
    fabric_llpp3_arprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp3_arqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp3_arsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp3_arvalid_s_o	: out std_logic := '0';
    fabric_llpp3_awaddr_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp3_awburst_s_o	: out std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp3_awcache_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp3_awid_s_o	: out std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp3_awlen_s_o	: out std_logic_vector(7   downto 0) := (others => '0');
    fabric_llpp3_awlock_s_o	: out std_logic := '0';
    fabric_llpp3_awprot_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp3_awqos_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp3_awsize_s_o	: out std_logic_vector(2   downto 0) := (others => '0');
    fabric_llpp3_awvalid_s_o	: out std_logic := '0';
    fabric_llpp3_bready_s_o	: out std_logic := '0';
    fabric_llpp3_rready_s_o	: out std_logic := '0';
    fabric_llpp3_wdata_s_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp3_wlast_s_o	: out std_logic := '0';
    fabric_llpp3_wstrb_s_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_llpp3_wvalid_s_o	: out std_logic := '0';
    fabric_llpp3_arready_s_i	: in std_logic := '0';
    fabric_llpp3_awready_s_i	: in std_logic := '0';
    fabric_llpp3_bid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp3_bresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp3_bvalid_s_i	: in std_logic := '0';
    fabric_llpp3_rdata_s_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_llpp3_rid_s_i	: in std_logic_vector(11  downto 0) := (others => '0');
    fabric_llpp3_rlast_s_i	: in std_logic := '0';
    fabric_llpp3_rresp_s_i	: in std_logic_vector(1   downto 0) := (others => '0');
    fabric_llpp3_rvalid_s_i	: in std_logic := '0';
    fabric_llpp3_wready_s_i	: in std_logic := '0';
    fabric_qos_pprdata_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_qos_ppready_o	: out std_logic := '0';
    fabric_qos_ppslverr_o	: out std_logic := '0';
    fabric_qos_pclk_i	: in std_logic := '0';
    fabric_qos_ppaddr_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_qos_ppenable_i	: in std_logic := '0';
    fabric_qos_ppwdata_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_qos_ppwrite_i	: in std_logic := '0';
    fabric_qos_presetn_i	: in std_logic := '0';
    fabric_qos_psel_i	: in std_logic := '0';
    fabric_tnd_hssl_flushin_o	: out std_logic := '0';
    fabric_tnd_hssl_trigin_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_paddr_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_fpga_apb_master_penable_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_psel_o	: out std_logic := '0';
    fabric_tnd_fpga_apb_master_pwdata_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_fpga_apb_master_pwrite_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_afvalid_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_atready_o	: out std_logic := '0';
    fabric_tnd_fpga_atb_master_syncreq_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_paddr_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_hssl_apb_master_penable_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_psel_o	: out std_logic := '0';
    fabric_tnd_hssl_apb_master_pwdata_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_hssl_apb_master_pwrite_o	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_afready_o	: out std_logic := '0';
    fabric_tnd_hssl_atb_master_atbytes_o	: out std_logic_vector(3   downto 0) := (others => '0');
    fabric_tnd_hssl_atb_master_atdata_o	: out std_logic_vector(127 downto 0) := (others => '0');
    fabric_tnd_hssl_atb_master_atid_o	: out std_logic_vector(6   downto 0) := (others => '0');
    fabric_tnd_hssl_atb_master_atvalid_o	: out std_logic := '0';
    fabric_tnd_trace_clk_traceoutportintf_o	: out std_logic := '0';
    fabric_tnd_trace_ctl_traceoutportintf_o	: out std_logic := '0';
    fabric_tnd_trace_data_traceoutportintf_o	: out std_logic_vector(31  downto 0) := (others => '0');
    fabric_tsvalue_tsgen_fpga_o	: out std_logic_vector(63  downto 0) := (others => '0');
    fabric_tnd_fpga_apb_master_prdata_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_fpga_apb_master_pready_i	: in std_logic := '0';
    fabric_tnd_fpga_apb_master_pslverr_i	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_afready_i	: in std_logic := '0';
    fabric_tnd_fpga_atb_master_atbytes_i	: in std_logic_vector(3   downto 0) := (others => '0');
    fabric_tnd_fpga_atb_master_atdata_i	: in std_logic_vector(127 downto 0) := (others => '0');
    fabric_tnd_fpga_atb_master_atid_i	: in std_logic_vector(6   downto 0) := (others => '0');
    fabric_tnd_fpga_atb_master_atvalid_i	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_prdata_i	: in std_logic_vector(31  downto 0) := (others => '0');
    fabric_tnd_hssl_apb_master_pready_i	: in std_logic := '0';
    fabric_tnd_hssl_apb_master_pslverr_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_afvalid_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_atready_i	: in std_logic := '0';
    fabric_tnd_hssl_atb_master_syncreq_i	: in std_logic := '0';
    fabric_watchdog0_signal_0_o	: out std_logic := '0';
    fabric_watchdog0_signal_1_o	: out std_logic := '0';
    fabric_watchdog1_signal_0_o	: out std_logic := '0';
    fabric_watchdog1_signal_1_o	: out std_logic := '0';
    fabric_watchdog2_signal_0_o	: out std_logic := '0';
    fabric_watchdog2_signal_1_o	: out std_logic := '0';
    fabric_watchdog3_signal_0_o	: out std_logic := '0';
    fabric_watchdog3_signal_1_o	: out std_logic := '0';
    fabric_tst_pll_lock_o	: out std_logic_vector(6   downto 0) := (others => '0');
    fabric_soc_mon_sensor_alarm_o	: out std_logic := '0';
    fabric_erom_fpga_cpu0_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu0_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu1_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu2_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_hiden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_hniden_i	: in std_logic := '0';
    fabric_erom_fpga_cpu3_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cs_dbgen_i	: in std_logic := '0';
    fabric_erom_fpga_cs_niden_i	: in std_logic := '0';
    fabric_erom_fpga_cs_deviceen_i	: in std_logic := '0';
    fabric_erom_fpga_cs_rst_n_i	: in std_logic := '0';
    fabric_erom_fpga_debug_en_i	: in std_logic := '0';
    fabric_enable_TMR_i	: in std_logic_vector(3   downto 0) := (others => '0')
);
end component NX_SOC_INTERFACE_WRAP;

component NX_BD is
generic (
    mode : string := "local_lowskew"
);
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_BD;

component NX_CY is
generic (
    add_carry  : integer := 0      -- 0: low - 1: high - 2: propagate
);
port (
    A1	: in std_logic := '0';
    A2	: in std_logic := '0';
    A3	: in std_logic := '0';
    A4	: in std_logic := '0';
    B1	: in std_logic := '0';
    B2	: in std_logic := '0';
    B3	: in std_logic := '0';
    B4	: in std_logic := '0';
    CI	: in std_logic := '0';
    CO	: out std_logic := '0';
    S1	: out std_logic := '0';
    S2	: out std_logic := '0';
    S3	: out std_logic := '0';
    S4	: out std_logic := '0'
);
end component NX_CY;

component NX_ECC is
port (
    CKD	: in std_logic := '0';
    CHK	: in std_logic := '0';
    COR	: out std_logic := '0';
    ERR	: out std_logic := '0'
    );
end component NX_ECC;

component NX_LUT is
generic (
    lut_table : bit_vector(15 downto 0) := B"0000000000000000" -- truthTable t15 ... t0
);
port (
    I1	: in std_logic := '0';
    I2	: in std_logic := '0';
    I3	: in std_logic := '0';
    I4	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_LUT;

component NX_DFF is
generic (
    dff_edge   : bit       := '0';
    dff_init   : bit       := '0';
    dff_load   : bit       := '0';
    dff_sync   : bit       := '0';
    dff_type   : integer   := 0;
    dff_ctxt   : std_logic := 'U'
);
port (
    I	: in std_logic := '0';
    CK	: in std_logic := '0';
    L	: in std_logic := '0';
    R	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_DFF;

component NX_BFF is
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_BFF;

component NX_DFR is
generic (
    location   : string  := "";
    iobname    : string  := "";
    path       : integer := 0;
    mode       : integer := 0;
    ring       : integer := 0;
    dff_edge   : bit     := '0';
    dff_init   : bit     := '0';
    dff_load   : bit     := '0';
    dff_sync   : bit     := '0';
    dff_type   : integer := 0
);
port (
    I	: in std_logic := '0';
    CK	: in std_logic := '0';
    L	: in std_logic := '0';
    R	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_DFR;

component NX_BFR is
generic (
    location   : string := "";
    iobname    : string := "";
    path       : integer := 0;
    mode       : integer := 0;
    data_inv   : bit     := '0';
    ring       : integer := 0
);
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_BFR;

component NX_IOB_I is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  1;
    locked               : bit     := '0'
);
port (
--  I  : in  std_logic;			// To prevent error in instanciation
    C	: in std_logic := '0';
    T	: in std_logic := '0';
    IO	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_IOB_I;

component NX_IOB_O is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  2;
    locked               : bit     := '0'
);
port (
    I	: in std_logic := '0';
    C	: in std_logic := '0';
    T	: in std_logic := '0';
--  O  : out std_logic;			// To prevent error in instanciation
    IO	: out std_logic := '0'
);
end component NX_IOB_O;

component NX_IOB is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  3;
    locked               : bit     := '0'
);
port (
    I	: in std_logic := '0';
    C	: in std_logic := '0';
    T	: in std_logic := '0';
    O	: out std_logic := '0';
    IO	: inout std_logic := '0'
);
end component NX_IOB;

-- beware following components are only intended for internal use. Do not try to instantiate them.
component NX_BUFFER is
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_BUFFER;

component NX_CSC is
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_CSC;

component NX_SCC is
port (
    I	: in std_logic := '0';
    O	: out std_logic := '0'
);
end component NX_SCC;

component NX_syn_tp is
port (
    I	: in std_logic := '0'
);
end component NX_syn_tp;

component NX_RAM is
generic (
   std_mode     : string := ""; -- standard mode [FAST_2kx18, SLOW_2kx18, NOECNOECC24, ...] empty for raw
   mcka_edge    : bit := '0';   -- 0: rising edge for port A clock - 1: falling edge
   mckb_edge    : bit := '0';   -- 0: rising edge for port B clock - 1: falling edge
   pcka_edge    : bit := '0';   -- 0: rising edge for pipe A clock - 1: falling edge
   pckb_edge    : bit := '0';   -- 0: rising edge for pipe B clock - 1: falling edge
   pipe_ia      : bit := '0';   -- 0: no pipe on port A input  - 1: pipe on port A input
   pipe_ib      : bit := '0';   -- 0: no pipe on port B input  - 1: pipe on port B input
   pipe_oa      : bit := '0';   -- 0: no pipe on port A output - 1: pipe on port A output
   pipe_ob      : bit := '0';   -- 0: no pipe on port B output - 1: pipe on port B output

   raw_config0  : bit_vector( 3 downto 0) := B"0000";			-- PRC
   raw_config1  : bit_vector(15 downto 0) := B"0000000000000000";	-- MOD

   -- For specific NG_LARGE Extended Features
   raw_l_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-LARGE extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_l_extend : bit_vector( 3 downto 0) := B"0000";	    -- Extended modes for NG-LARGE (Scrubbing, test... )

   -- For specific NG_ULTRA Extended Features
   raw_u_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-ULTRA extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_u_extend : bit_vector( 7 downto 0) := B"00000000";   -- Extended modes for NG-ULTRA (Scrubbing, test... )

   mem_ctxt     : string := ""				    -- context initialization
   );
port (
    ACK	: in std_logic := '0';
    ACKC	: in std_logic := '0';
    ACKD	: in std_logic := '0';
    ACKR	: in std_logic := '0';
    BCK	: in std_logic := '0';
    BCKC	: in std_logic := '0';
    BCKD	: in std_logic := '0';
    BCKR	: in std_logic := '0';

    AI1	: in std_logic := '0';
    AI2	: in std_logic := '0';
    AI3	: in std_logic := '0';
    AI4	: in std_logic := '0';
    AI5	: in std_logic := '0';
    AI6	: in std_logic := '0';
    AI7	: in std_logic := '0';
    AI8	: in std_logic := '0';
    AI9	: in std_logic := '0';
    AI10	: in std_logic := '0';
    AI11	: in std_logic := '0';
    AI12	: in std_logic := '0';
    AI13	: in std_logic := '0';
    AI14	: in std_logic := '0';
    AI15	: in std_logic := '0';
    AI16	: in std_logic := '0';

    AI17	: in std_logic := '0';
    AI18	: in std_logic := '0';
    AI19	: in std_logic := '0';
    AI20	: in std_logic := '0';
    AI21	: in std_logic := '0';
    AI22	: in std_logic := '0';
    AI23	: in std_logic := '0';
    AI24	: in std_logic := '0';

    BI1	: in std_logic := '0';
    BI2	: in std_logic := '0';
    BI3	: in std_logic := '0';
    BI4	: in std_logic := '0';
    BI5	: in std_logic := '0';
    BI6	: in std_logic := '0';
    BI7	: in std_logic := '0';
    BI8	: in std_logic := '0';
    BI9	: in std_logic := '0';
    BI10	: in std_logic := '0';
    BI11	: in std_logic := '0';
    BI12	: in std_logic := '0';
    BI13	: in std_logic := '0';
    BI14	: in std_logic := '0';
    BI15	: in std_logic := '0';
    BI16	: in std_logic := '0';

    BI17	: in std_logic := '0';
    BI18	: in std_logic := '0';
    BI19	: in std_logic := '0';
    BI20	: in std_logic := '0';
    BI21	: in std_logic := '0';
    BI22	: in std_logic := '0';
    BI23	: in std_logic := '0';
    BI24	: in std_logic := '0';

    ACOR	: out std_logic := '0';
    AERR	: out std_logic := '0';
    BCOR	: out std_logic := '0';
    BERR	: out std_logic := '0';

    AO1	: out std_logic := '0';
    AO2	: out std_logic := '0';
    AO3	: out std_logic := '0';
    AO4	: out std_logic := '0';
    AO5	: out std_logic := '0';
    AO6	: out std_logic := '0';
    AO7	: out std_logic := '0';
    AO8	: out std_logic := '0';
    AO9	: out std_logic := '0';
    AO10	: out std_logic := '0';
    AO11	: out std_logic := '0';
    AO12	: out std_logic := '0';
    AO13	: out std_logic := '0';
    AO14	: out std_logic := '0';
    AO15	: out std_logic := '0';
    AO16	: out std_logic := '0';

    AO17	: out std_logic := '0';
    AO18	: out std_logic := '0';
    AO19	: out std_logic := '0';
    AO20	: out std_logic := '0';
    AO21	: out std_logic := '0';
    AO22	: out std_logic := '0';
    AO23	: out std_logic := '0';
    AO24	: out std_logic := '0';

    BO1	: out std_logic := '0';
    BO2	: out std_logic := '0';
    BO3	: out std_logic := '0';
    BO4	: out std_logic := '0';
    BO5	: out std_logic := '0';
    BO6	: out std_logic := '0';
    BO7	: out std_logic := '0';
    BO8	: out std_logic := '0';
    BO9	: out std_logic := '0';
    BO10	: out std_logic := '0';
    BO11	: out std_logic := '0';
    BO12	: out std_logic := '0';
    BO13	: out std_logic := '0';
    BO14	: out std_logic := '0';
    BO15	: out std_logic := '0';
    BO16	: out std_logic := '0';

    BO17	: out std_logic := '0';
    BO18	: out std_logic := '0';
    BO19	: out std_logic := '0';
    BO20	: out std_logic := '0';
    BO21	: out std_logic := '0';
    BO22	: out std_logic := '0';
    BO23	: out std_logic := '0';
    BO24	: out std_logic := '0';

    AA1	: in std_logic := '0';
    AA2	: in std_logic := '0';
    AA3	: in std_logic := '0';
    AA4	: in std_logic := '0';
    AA5	: in std_logic := '0';
    AA6	: in std_logic := '0';

    AA7	: in std_logic := '0';
    AA8	: in std_logic := '0';
    AA9	: in std_logic := '0';
    AA10	: in std_logic := '0';
    AA11	: in std_logic := '0';
    AA12	: in std_logic := '0';
    AA13	: in std_logic := '0';
    AA14	: in std_logic := '0';
    AA15	: in std_logic := '0';
    AA16	: in std_logic := '0';

    ACS	: in std_logic := '0';
    AWE	: in std_logic := '0';
    AR	: in std_logic := '0';

    BA1	: in std_logic := '0';
    BA2	: in std_logic := '0';
    BA3	: in std_logic := '0';
    BA4	: in std_logic := '0';
    BA5	: in std_logic := '0';
    BA6	: in std_logic := '0';

    BA7	: in std_logic := '0';
    BA8	: in std_logic := '0';
    BA9	: in std_logic := '0';
    BA10	: in std_logic := '0';
    BA11	: in std_logic := '0';
    BA12	: in std_logic := '0';
    BA13	: in std_logic := '0';
    BA14	: in std_logic := '0';
    BA15	: in std_logic := '0';
    BA16	: in std_logic := '0';

    BCS	: in std_logic := '0';
    BWE	: in std_logic := '0';
    BR	: in std_logic := '0'
);
end component NX_RAM;

component NX_RAM_WRAP is
generic (
   std_mode     : string := ""; -- standard mode [FAST_2kx18, SLOW_2kx18, NOECNOECC24, ...] empty for raw
   mcka_edge    : bit := '0';   -- 0: rising edge for port A clock - 1: falling edge
   mckb_edge    : bit := '0';   -- 0: rising edge for port B clock - 1: falling edge
   pcka_edge    : bit := '0';   -- 0: rising edge for pipe A clock - 1: falling edge
   pckb_edge    : bit := '0';   -- 0: rising edge for pipe B clock - 1: falling edge

   pipe_ia      : bit := '0';   -- 0: no pipe on port A input  - 1: pipe on port A input
   pipe_ib      : bit := '0';   -- 0: no pipe on port B input  - 1: pipe on port B input
   pipe_oa      : bit := '0';   -- 0: no pipe on port A output - 1: pipe on port A output
   pipe_ob      : bit := '0';   -- 0: no pipe on port B output - 1: pipe on port B output

   raw_config0  : bit_vector( 3 downto 0) := B"0000";			-- PRC
   raw_config1  : bit_vector(15 downto 0) := B"0000000000000000";	-- MOD

   -- For specific NG_LARGE Extended Features
   raw_l_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-LARGE extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_l_extend : bit_vector( 3 downto 0) := B"0000";	    -- Extended modes for NG-LARGE (Scrubbing, test... )

   -- For specific NG_ULTRA Extended Features
   raw_u_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-ULTRA extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_u_extend : bit_vector( 7 downto 0) := B"00000000";   -- Extended modes for NG-ULTRA (Scrubbing, test... )

   mem_ctxt     : string := ""				    -- context initialization
);
port (
    ACK	: in std_logic := '0';
    ACKD	: in std_logic := '0';
    ACKR	: in std_logic := '0';
    BCK	: in std_logic := '0';
    BCKD	: in std_logic := '0';
    BCKR	: in std_logic := '0';

    AI	: in std_logic_vector(23 downto 0) := (others => '0');
    BI	: in std_logic_vector(23 downto 0) := (others => '0');

    ACOR	: out std_logic := '0';
    AERR	: out std_logic := '0';
    BCOR	: out std_logic := '0';
    BERR	: out std_logic := '0';

    AO	: out std_logic_vector(23 downto 0) := (others => '0');
    BO	: out std_logic_vector(23 downto 0) := (others => '0');
    AA	: in std_logic_vector(15 downto 0) := (others => '0');

    ACS	: in std_logic := '0';
    AWE	: in std_logic := '0';
    AR	: in std_logic := '0';

    BA	: in std_logic_vector(15 downto 0) := (others => '0');

    BCS	: in std_logic := '0';
    BWE	: in std_logic := '0';
    BR	: in std_logic := '0'
);
end component NX_RAM_WRAP;


end nxPackage;
-- =================================================================================================
--   NX_CDC_L definition                                                                2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CDC_L is
generic (
    mode : bit := '0';
    rck_edge : bit := '0';
    wck_edge : bit := '0'
);
port (
    CK  : in  std_logic;
    RI1 : in  std_logic;
    RI2 : in  std_logic;
    RI3 : in  std_logic;
    RI4 : in  std_logic;
    RI5 : in  std_logic;
    RI6 : in  std_logic;
    RO1 : out std_logic;
    RO2 : out std_logic;
    RO3 : out std_logic;
    RO4 : out std_logic;
    RO5 : out std_logic;
    RO6 : out std_logic;
    WI1 : in  std_logic;
    WI2 : in  std_logic;
    WI3 : in  std_logic;
    WI4 : in  std_logic;
    WI5 : in  std_logic;
    WI6 : in  std_logic;
    WO1 : out std_logic;
    WO2 : out std_logic;
    WO3 : out std_logic;
    WO4 : out std_logic;
    WO5 : out std_logic;
    WO6 : out std_logic
);
end NX_CDC_L;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_FIFO_CDC_L definition                                                           2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_FIFO_CDC_L is
generic (
    mode : bit := '1'
);
port (
    XRCK : in  std_logic;
    XWCK : in  std_logic;
    XRI1 : in  std_logic;
    XRI2 : in  std_logic;
    XRI3 : in  std_logic;
    XRI4 : in  std_logic;
    XRI5 : in  std_logic;
    XRI6 : in  std_logic;
    XWI1 : in  std_logic;
    XWI2 : in  std_logic;
    XWI3 : in  std_logic;
    XWI4 : in  std_logic;
    XWI5 : in  std_logic;
    XWI6 : in  std_logic;
    RO1  : out std_logic;
    RO2  : out std_logic;
    RO3  : out std_logic;
    RO4  : out std_logic;
    RO5  : out std_logic;
    RO6  : out std_logic;
    WO1  : out std_logic;
    WO2  : out std_logic;
    WO3  : out std_logic;
    WO4  : out std_logic;
    WO5  : out std_logic;
    WO6  : out std_logic
);
end NX_FIFO_CDC_L;
-- =================================================================================================
--   NX_DSPDPRAM_FULL_L definition                                                       2020/02/03
-- =================================================================================================

-- NX_DSPDPRAM_FULL_L#{{{#
library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DSPDPRAM_FULL_L is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    dsp0_clk_i  : in  std_logic;                                        -- DSP1.CK
    dsp0_rst_i  : in  std_logic; -- rst_i  et rstsys_i                  -- DSP1.R
    dsp0_rstz_i : in  std_logic; -- rstz_i et rstzsys_i                 -- DSP1.RZ
    dsp0_we_i   : in  std_logic; -- we_i   et wesys_i                   -- DSP1.WE
    dsp0_cy_i   : in  std_logic;                                        -- DSP1.CI
    dsp0_a_i    : in  std_logic_vector(23 downto 0);                    -- DSP1.A
    dsp0_b_i    : in  std_logic_vector(17 downto 0);                    -- DSP1.B
    dsp0_c_i    : in  std_logic_vector(35 downto 0);                    -- DSP1.C
    dsp0_d_i    : in  std_logic_vector(17 downto 0);                    -- DSP1.D

    dsp0_z_o    : out std_logic_vector(55 downto 0);                    -- DSP1.Z
    dsp0_cy_o   : out std_logic;                                        -- DSP1.CO
    dsp0_cy36_o : out std_logic;                                        -- DSP1.CO37
    dsp0_cy56_o : out std_logic;                                        -- DSP1.CO57
    dsp0_ovf_o  : out std_logic;                                        -- DSP1.OVF

    dsp1_clk_i  : in  std_logic;                                        -- DSP2.CK
    dsp1_rst_i  : in  std_logic; -- rst_i  et rstsys_i                  -- DSP2.R
    dsp1_rstz_i : in  std_logic; -- rstz_i et rstzsys_i                 -- DSP2.RZ
    dsp1_we_i   : in  std_logic; -- we_i   et wesys_i                   -- DSP2.WE
    dsp1_cy_i   : in  std_logic;                                        -- DSP2.CI
    dsp1_a_i    : in  std_logic_vector(23 downto 0);                    -- DSP2.A
    dsp1_b_i    : in  std_logic_vector(17 downto 0);                    -- DSP2.B
    dsp1_c_i    : in  std_logic_vector(35 downto 0);                    -- DSP2.C
    dsp1_d_i    : in  std_logic_vector(17 downto 0);                    -- DSP2.D

    dsp1_z_o    : out std_logic_vector(55 downto 0);                    -- DSP2.Z
    dsp1_cy_o   : out std_logic;                                        -- DSP2.CO
    dsp1_cy36_o : out std_logic;                                        -- DSP2.CO37
    dsp1_cy56_o : out std_logic;                                        -- DSP2.CO57
    dsp1_ovf_o  : out std_logic;                                        -- DSP2.OVF

    dsp_ca_i    : in  std_logic_vector(23 downto 0);                    -- DSP2.CAI
    dsp_cb_i    : in  std_logic_vector(17 downto 0);                    -- DSP2.CBI
    dsp_cz_i    : in  std_logic_vector(55 downto 0);                    -- DSP2.CZI
    dsp_ccy_i   : in  std_logic;                                        -- DSP1.CCI
    dsp_ca_o    : out std_logic_vector(23 downto 0);                    -- DSP1.CAO
    dsp_cb_o    : out std_logic_vector(17 downto 0);                    -- DSP1.CBO
    dsp_cz_o    : out std_logic_vector(55 downto 0);                    -- DSP1.CZO
    dsp_ccy_o   : out std_logic;                                        -- DSP2.CCO


    dpram_clkmem0_i          : in  std_logic;                           -- RAM.ACK
    dpram_clkmemclone0_i     : in  std_logic;                           -- RAM.ACKC
    dpram_clkmem90_0_i       : in  std_logic;                           -- RAM.ACKD
    dpram_clkreg0_i          : in  std_logic;                           -- RAM.ACKR
    dpram_rst0_i             : in  std_logic; -- rst_i et rstsys_i      -- RAM.AR
    dpram_cs0_i              : in  std_logic; -- cs_i  et cssys_i       -- RAM.ACS
    dpram_we0_i              : in  std_logic; -- we_i  et wesys_i       -- RAM.AWE
    dpram_addr0_i            : in  std_logic_vector(15 downto 0);       -- RAM.AA
    dpram_din0_i             : in  std_logic_vector(23 downto 0);       -- RAM.AI
    dpram_dout0_o            : out std_logic_vector(23 downto 0);       -- RAM.AO
    dpram_ecc_corrected0_o   : out std_logic;                           -- RAM.ACOR
    dpram_ecc_uncorrected0_o : out std_logic;                           -- RAM.AERR

    dpram_clkmem1_i          : in  std_logic;                           -- RAM.BCK
    dpram_clkmemclone1_i     : in  std_logic;                           -- RAM.BCKC
    dpram_clkmem90_1_i       : in  std_logic;                           -- RAM.BCKD
    dpram_clkreg1_i          : in  std_logic;                           -- RAM.BCKR
    dpram_rst1_i             : in  std_logic; -- rst_i et rstsys_i      -- RAM.BR
    dpram_cs1_i              : in  std_logic; -- cs_i  et cssys_i       -- RAM.BCS
    dpram_we1_i              : in  std_logic; -- we_i  et wesys_i       -- RAM.BWE
    dpram_addr1_i            : in  std_logic_vector(15 downto 0);       -- RAM.BA
    dpram_din1_i             : in  std_logic_vector(23 downto 0);       -- RAM.BI
    dpram_dout1_o            : out std_logic_vector(23 downto 0);       -- RAM.BO
    dpram_ecc_corrected1_o   : out std_logic;                           -- RAM.BCOR
    dpram_ecc_uncorrected1_o : out std_logic                            -- RAM.BERR
);
end NX_DSPDPRAM_FULL_L;
--#}}}#

-- architecture NX_RTL of NX_DSPDPRAM_FULL_L#{{{#
architecture NX_RTL of NX_DSPDPRAM_FULL_L is

  -- component NX_DSP_L_BOX#{{{#
  component NX_DSP_L_BOX
  generic (
      col    : integer := 2;
      row    : integer := 4;
      cfg0_i : bit_vector(95 downto 0) := (others => '0');
      cfg1_i : bit_vector(95 downto 0) := (others => '0')
  );
  port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
  );
  end component;
  --#}}}#

  -- component NX_RAM_L_BOX#{{{#
  component NX_RAM_L_BOX
  generic (
      col    : integer := 2;
      row    : integer := 4;
      cfg0_i : bit_vector(95 downto 0) := (others => '0');
      cfg1_i : bit_vector(95 downto 0) := (others => '0')
  );
  port (
    ACK   : in  std_logic;
    ACKC  : in  std_logic;
    ACKD  : in  std_logic;
    ACKR  : in  std_logic;
    BCK   : in  std_logic;
    BCKC  : in  std_logic;
    BCKD  : in  std_logic;
    BCKR  : in  std_logic;

    AI1   : in  std_logic;
    AI2   : in  std_logic;
    AI3   : in  std_logic;
    AI4   : in  std_logic;
    AI5   : in  std_logic;
    AI6   : in  std_logic;
    AI7   : in  std_logic;
    AI8   : in  std_logic;
    AI9   : in  std_logic;
    AI10  : in  std_logic;
    AI11  : in  std_logic;
    AI12  : in  std_logic;
    AI13  : in  std_logic;
    AI14  : in  std_logic;
    AI15  : in  std_logic;
    AI16  : in  std_logic;

    AI17  : in  std_logic;
    AI18  : in  std_logic;
    AI19  : in  std_logic;
    AI20  : in  std_logic;
    AI21  : in  std_logic;
    AI22  : in  std_logic;
    AI23  : in  std_logic;
    AI24  : in  std_logic;

    BI1   : in  std_logic;
    BI2   : in  std_logic;
    BI3   : in  std_logic;
    BI4   : in  std_logic;
    BI5   : in  std_logic;
    BI6   : in  std_logic;
    BI7   : in  std_logic;
    BI8   : in  std_logic;
    BI9   : in  std_logic;
    BI10  : in  std_logic;
    BI11  : in  std_logic;
    BI12  : in  std_logic;
    BI13  : in  std_logic;
    BI14  : in  std_logic;
    BI15  : in  std_logic;
    BI16  : in  std_logic;

    BI17  : in  std_logic;
    BI18  : in  std_logic;
    BI19  : in  std_logic;
    BI20  : in  std_logic;
    BI21  : in  std_logic;
    BI22  : in  std_logic;
    BI23  : in  std_logic;
    BI24  : in  std_logic;

    ACOR  : out std_logic;
    AERR  : out std_logic;
    BCOR  : out std_logic;
    BERR  : out std_logic;

    AO1   : out std_logic;
    AO2   : out std_logic;
    AO3   : out std_logic;
    AO4   : out std_logic;
    AO5   : out std_logic;
    AO6   : out std_logic;
    AO7   : out std_logic;
    AO8   : out std_logic;
    AO9   : out std_logic;
    AO10  : out std_logic;
    AO11  : out std_logic;
    AO12  : out std_logic;
    AO13  : out std_logic;
    AO14  : out std_logic;
    AO15  : out std_logic;
    AO16  : out std_logic;

    AO17  : out std_logic;
    AO18  : out std_logic;
    AO19  : out std_logic;
    AO20  : out std_logic;
    AO21  : out std_logic;
    AO22  : out std_logic;
    AO23  : out std_logic;
    AO24  : out std_logic;

    BO1   : out std_logic;
    BO2   : out std_logic;
    BO3   : out std_logic;
    BO4   : out std_logic;
    BO5   : out std_logic;
    BO6   : out std_logic;
    BO7   : out std_logic;
    BO8   : out std_logic;
    BO9   : out std_logic;
    BO10  : out std_logic;
    BO11  : out std_logic;
    BO12  : out std_logic;
    BO13  : out std_logic;
    BO14  : out std_logic;
    BO15  : out std_logic;
    BO16  : out std_logic;

    BO17  : out std_logic;
    BO18  : out std_logic;
    BO19  : out std_logic;
    BO20  : out std_logic;
    BO21  : out std_logic;
    BO22  : out std_logic;
    BO23  : out std_logic;
    BO24  : out std_logic;

    AA1   : in  std_logic;
    AA2   : in  std_logic;
    AA3   : in  std_logic;
    AA4   : in  std_logic;
    AA5   : in  std_logic;
    AA6   : in  std_logic;

    AA7   : in  std_logic;
    AA8   : in  std_logic;
    AA9   : in  std_logic;
    AA10  : in  std_logic;
    AA11  : in  std_logic;
    AA12  : in  std_logic;
    AA13  : in  std_logic;
    AA14  : in  std_logic;
    AA15  : in  std_logic;
    AA16  : in  std_logic;

    ACS   : in  std_logic;
    AWE   : in  std_logic;
    AR    : in  std_logic;

    BA1   : in  std_logic;
    BA2   : in  std_logic;
    BA3   : in  std_logic;
    BA4   : in  std_logic;
    BA5   : in  std_logic;
    BA6   : in  std_logic;

    BA7   : in  std_logic;
    BA8   : in  std_logic;
    BA9   : in  std_logic;
    BA10  : in  std_logic;
    BA11  : in  std_logic;
    BA12  : in  std_logic;
    BA13  : in  std_logic;
    BA14  : in  std_logic;
    BA15  : in  std_logic;
    BA16  : in  std_logic;

    BCS   : in  std_logic;
    BWE   : in  std_logic;
    BR    : in  std_logic
  );
  end component;
  --#}}}#

signal c_cy_int : std_logic;
signal c_a_int : std_logic_vector(23 downto 0);
signal c_b_int : std_logic_vector(17 downto 0);
signal c_z_int : std_logic_vector(55 downto 0);

attribute syn_preserve : boolean;
attribute syn_preserve of dsp_0 : label is true;
attribute syn_preserve of dsp_1 : label is true;
attribute syn_preserve of ram_0 : label is true;

begin

-- instance dsp0#{{{#
dsp_0 : NX_DSP_L_BOX
generic map (
    col    => col
  , row    => row
  , cfg0_i => cfg0_i
  , cfg1_i => cfg1_i
)
port map (
      A1    => dsp0_a_i(0)
   ,  A2    => dsp0_a_i(1)
   ,  A3    => dsp0_a_i(2)
   ,  A4    => dsp0_a_i(3)
   ,  A5    => dsp0_a_i(4)
   ,  A6    => dsp0_a_i(5)
   ,  A7    => dsp0_a_i(6)
   ,  A8    => dsp0_a_i(7)
   ,  A9    => dsp0_a_i(8)
   ,  A10   => dsp0_a_i(9)
   ,  A11   => dsp0_a_i(10)
   ,  A12   => dsp0_a_i(11)
   ,  A13   => dsp0_a_i(12)
   ,  A14   => dsp0_a_i(13)
   ,  A15   => dsp0_a_i(14)
   ,  A16   => dsp0_a_i(15)
   ,  A17   => dsp0_a_i(16)
   ,  A18   => dsp0_a_i(17)
   ,  A19   => dsp0_a_i(18)
   ,  A20   => dsp0_a_i(19)
   ,  A21   => dsp0_a_i(20)
   ,  A22   => dsp0_a_i(21)
   ,  A23   => dsp0_a_i(22)
   ,  A24   => dsp0_a_i(23)
   ,  B1    => dsp0_b_i(0)
   ,  B2    => dsp0_b_i(1)
   ,  B3    => dsp0_b_i(2)
   ,  B4    => dsp0_b_i(3)
   ,  B5    => dsp0_b_i(4)
   ,  B6    => dsp0_b_i(5)
   ,  B7    => dsp0_b_i(6)
   ,  B8    => dsp0_b_i(7)
   ,  B9    => dsp0_b_i(8)
   ,  B10   => dsp0_b_i(9)
   ,  B11   => dsp0_b_i(10)
   ,  B12   => dsp0_b_i(11)
   ,  B13   => dsp0_b_i(12)
   ,  B14   => dsp0_b_i(13)
   ,  B15   => dsp0_b_i(14)
   ,  B16   => dsp0_b_i(15)
   ,  B17   => dsp0_b_i(16)
   ,  B18   => dsp0_b_i(17)
   ,  C1    => dsp0_c_i(0)
   ,  C2    => dsp0_c_i(1)
   ,  C3    => dsp0_c_i(2)
   ,  C4    => dsp0_c_i(3)
   ,  C5    => dsp0_c_i(4)
   ,  C6    => dsp0_c_i(5)
   ,  C7    => dsp0_c_i(6)
   ,  C8    => dsp0_c_i(7)
   ,  C9    => dsp0_c_i(8)
   ,  C10   => dsp0_c_i(9)
   ,  C11   => dsp0_c_i(10)
   ,  C12   => dsp0_c_i(11)
   ,  C13   => dsp0_c_i(12)
   ,  C14   => dsp0_c_i(13)
   ,  C15   => dsp0_c_i(14)
   ,  C16   => dsp0_c_i(15)
   ,  C17   => dsp0_c_i(16)
   ,  C18   => dsp0_c_i(17)
   ,  C19   => dsp0_c_i(18)
   ,  C20   => dsp0_c_i(19)
   ,  C21   => dsp0_c_i(20)
   ,  C22   => dsp0_c_i(21)
   ,  C23   => dsp0_c_i(22)
   ,  C24   => dsp0_c_i(23)
   ,  C25   => dsp0_c_i(24)
   ,  C26   => dsp0_c_i(25)
   ,  C27   => dsp0_c_i(26)
   ,  C28   => dsp0_c_i(27)
   ,  C29   => dsp0_c_i(28)
   ,  C30   => dsp0_c_i(29)
   ,  C31   => dsp0_c_i(30)
   ,  C32   => dsp0_c_i(31)
   ,  C33   => dsp0_c_i(32)
   ,  C34   => dsp0_c_i(33)
   ,  C35   => dsp0_c_i(34)
   ,  C36   => dsp0_c_i(35)
   ,  CAI1  => c_a_int(0)
   ,  CAI2  => c_a_int(1)
   ,  CAI3  => c_a_int(2)
   ,  CAI4  => c_a_int(3)
   ,  CAI5  => c_a_int(4)
   ,  CAI6  => c_a_int(5)
   ,  CAI7  => c_a_int(6)
   ,  CAI8  => c_a_int(7)
   ,  CAI9  => c_a_int(8)
   ,  CAI10 => c_a_int(9)
   ,  CAI11 => c_a_int(10)
   ,  CAI12 => c_a_int(11)
   ,  CAI13 => c_a_int(12)
   ,  CAI14 => c_a_int(13)
   ,  CAI15 => c_a_int(14)
   ,  CAI16 => c_a_int(15)
   ,  CAI17 => c_a_int(16)
   ,  CAI18 => c_a_int(17)
   ,  CAI19 => c_a_int(18)
   ,  CAI20 => c_a_int(19)
   ,  CAI21 => c_a_int(20)
   ,  CAI22 => c_a_int(21)
   ,  CAI23 => c_a_int(22)
   ,  CAI24 => c_a_int(23)
   ,  CAO1  => dsp_ca_o(0)
   ,  CAO2  => dsp_ca_o(1)
   ,  CAO3  => dsp_ca_o(2)
   ,  CAO4  => dsp_ca_o(3)
   ,  CAO5  => dsp_ca_o(4)
   ,  CAO6  => dsp_ca_o(5)
   ,  CAO7  => dsp_ca_o(6)
   ,  CAO8  => dsp_ca_o(7)
   ,  CAO9  => dsp_ca_o(8)
   ,  CAO10 => dsp_ca_o(9)
   ,  CAO11 => dsp_ca_o(10)
   ,  CAO12 => dsp_ca_o(11)
   ,  CAO13 => dsp_ca_o(12)
   ,  CAO14 => dsp_ca_o(13)
   ,  CAO15 => dsp_ca_o(14)
   ,  CAO16 => dsp_ca_o(15)
   ,  CAO17 => dsp_ca_o(16)
   ,  CAO18 => dsp_ca_o(17)
   ,  CAO19 => dsp_ca_o(18)
   ,  CAO20 => dsp_ca_o(19)
   ,  CAO21 => dsp_ca_o(20)
   ,  CAO22 => dsp_ca_o(21)
   ,  CAO23 => dsp_ca_o(22)
   ,  CAO24 => dsp_ca_o(23)
   ,  CBI1  => c_b_int(0)
   ,  CBI2  => c_b_int(1)
   ,  CBI3  => c_b_int(2)
   ,  CBI4  => c_b_int(3)
   ,  CBI5  => c_b_int(4)
   ,  CBI6  => c_b_int(5)
   ,  CBI7  => c_b_int(6)
   ,  CBI8  => c_b_int(7)
   ,  CBI9  => c_b_int(8)
   ,  CBI10 => c_b_int(9)
   ,  CBI11 => c_b_int(10)
   ,  CBI12 => c_b_int(11)
   ,  CBI13 => c_b_int(12)
   ,  CBI14 => c_b_int(13)
   ,  CBI15 => c_b_int(14)
   ,  CBI16 => c_b_int(15)
   ,  CBI17 => c_b_int(16)
   ,  CBI18 => c_b_int(17)
   ,  CBO1  => dsp_cb_o(0)
   ,  CBO2  => dsp_cb_o(1)
   ,  CBO3  => dsp_cb_o(2)
   ,  CBO4  => dsp_cb_o(3)
   ,  CBO5  => dsp_cb_o(4)
   ,  CBO6  => dsp_cb_o(5)
   ,  CBO7  => dsp_cb_o(6)
   ,  CBO8  => dsp_cb_o(7)
   ,  CBO9  => dsp_cb_o(8)
   ,  CBO10 => dsp_cb_o(9)
   ,  CBO11 => dsp_cb_o(10)
   ,  CBO12 => dsp_cb_o(11)
   ,  CBO13 => dsp_cb_o(12)
   ,  CBO14 => dsp_cb_o(13)
   ,  CBO15 => dsp_cb_o(14)
   ,  CBO16 => dsp_cb_o(15)
   ,  CBO17 => dsp_cb_o(16)
   ,  CBO18 => dsp_cb_o(17)
   ,  CCI   => dsp_ccy_i
   ,  CCO   => c_cy_int
   ,  CI    => dsp0_cy_i
   ,  CK    => dsp0_clk_i
   ,  CO    => dsp0_cy_o
   ,  CO37  => dsp0_cy36_o
   ,  CO57  => dsp0_cy56_o
   ,  CZI1  => c_z_int(0)
   ,  CZI2  => c_z_int(1)
   ,  CZI3  => c_z_int(2)
   ,  CZI4  => c_z_int(3)
   ,  CZI5  => c_z_int(4)
   ,  CZI6  => c_z_int(5)
   ,  CZI7  => c_z_int(6)
   ,  CZI8  => c_z_int(7)
   ,  CZI9  => c_z_int(8)
   ,  CZI10 => c_z_int(9)
   ,  CZI11 => c_z_int(10)
   ,  CZI12 => c_z_int(11)
   ,  CZI13 => c_z_int(12)
   ,  CZI14 => c_z_int(13)
   ,  CZI15 => c_z_int(14)
   ,  CZI16 => c_z_int(15)
   ,  CZI17 => c_z_int(16)
   ,  CZI18 => c_z_int(17)
   ,  CZI19 => c_z_int(18)
   ,  CZI20 => c_z_int(19)
   ,  CZI21 => c_z_int(20)
   ,  CZI22 => c_z_int(21)
   ,  CZI23 => c_z_int(22)
   ,  CZI24 => c_z_int(23)
   ,  CZI25 => c_z_int(24)
   ,  CZI26 => c_z_int(25)
   ,  CZI27 => c_z_int(26)
   ,  CZI28 => c_z_int(27)
   ,  CZI29 => c_z_int(28)
   ,  CZI30 => c_z_int(29)
   ,  CZI31 => c_z_int(30)
   ,  CZI32 => c_z_int(31)
   ,  CZI33 => c_z_int(32)
   ,  CZI34 => c_z_int(33)
   ,  CZI35 => c_z_int(34)
   ,  CZI36 => c_z_int(35)
   ,  CZI37 => c_z_int(36)
   ,  CZI38 => c_z_int(37)
   ,  CZI39 => c_z_int(38)
   ,  CZI40 => c_z_int(39)
   ,  CZI41 => c_z_int(40)
   ,  CZI42 => c_z_int(41)
   ,  CZI43 => c_z_int(42)
   ,  CZI44 => c_z_int(43)
   ,  CZI45 => c_z_int(44)
   ,  CZI46 => c_z_int(45)
   ,  CZI47 => c_z_int(46)
   ,  CZI48 => c_z_int(47)
   ,  CZI49 => c_z_int(48)
   ,  CZI50 => c_z_int(49)
   ,  CZI51 => c_z_int(50)
   ,  CZI52 => c_z_int(51)
   ,  CZI53 => c_z_int(52)
   ,  CZI54 => c_z_int(53)
   ,  CZI55 => c_z_int(54)
   ,  CZI56 => c_z_int(55)
   ,  CZO1  => dsp_cz_o(0)
   ,  CZO2  => dsp_cz_o(1)
   ,  CZO3  => dsp_cz_o(2)
   ,  CZO4  => dsp_cz_o(3)
   ,  CZO5  => dsp_cz_o(4)
   ,  CZO6  => dsp_cz_o(5)
   ,  CZO7  => dsp_cz_o(6)
   ,  CZO8  => dsp_cz_o(7)
   ,  CZO9  => dsp_cz_o(8)
   ,  CZO10 => dsp_cz_o(9)
   ,  CZO11 => dsp_cz_o(10)
   ,  CZO12 => dsp_cz_o(11)
   ,  CZO13 => dsp_cz_o(12)
   ,  CZO14 => dsp_cz_o(13)
   ,  CZO15 => dsp_cz_o(14)
   ,  CZO16 => dsp_cz_o(15)
   ,  CZO17 => dsp_cz_o(16)
   ,  CZO18 => dsp_cz_o(17)
   ,  CZO19 => dsp_cz_o(18)
   ,  CZO20 => dsp_cz_o(19)
   ,  CZO21 => dsp_cz_o(20)
   ,  CZO22 => dsp_cz_o(21)
   ,  CZO23 => dsp_cz_o(22)
   ,  CZO24 => dsp_cz_o(23)
   ,  CZO25 => dsp_cz_o(24)
   ,  CZO26 => dsp_cz_o(25)
   ,  CZO27 => dsp_cz_o(26)
   ,  CZO28 => dsp_cz_o(27)
   ,  CZO29 => dsp_cz_o(28)
   ,  CZO30 => dsp_cz_o(29)
   ,  CZO31 => dsp_cz_o(30)
   ,  CZO32 => dsp_cz_o(31)
   ,  CZO33 => dsp_cz_o(32)
   ,  CZO34 => dsp_cz_o(33)
   ,  CZO35 => dsp_cz_o(34)
   ,  CZO36 => dsp_cz_o(35)
   ,  CZO37 => dsp_cz_o(36)
   ,  CZO38 => dsp_cz_o(37)
   ,  CZO39 => dsp_cz_o(38)
   ,  CZO40 => dsp_cz_o(39)
   ,  CZO41 => dsp_cz_o(40)
   ,  CZO42 => dsp_cz_o(41)
   ,  CZO43 => dsp_cz_o(42)
   ,  CZO44 => dsp_cz_o(43)
   ,  CZO45 => dsp_cz_o(44)
   ,  CZO46 => dsp_cz_o(45)
   ,  CZO47 => dsp_cz_o(46)
   ,  CZO48 => dsp_cz_o(47)
   ,  CZO49 => dsp_cz_o(48)
   ,  CZO50 => dsp_cz_o(49)
   ,  CZO51 => dsp_cz_o(50)
   ,  CZO52 => dsp_cz_o(51)
   ,  CZO53 => dsp_cz_o(52)
   ,  CZO54 => dsp_cz_o(53)
   ,  CZO55 => dsp_cz_o(54)
   ,  CZO56 => dsp_cz_o(55)
   ,  D1    => dsp0_d_i(0)
   ,  D2    => dsp0_d_i(1)
   ,  D3    => dsp0_d_i(2)
   ,  D4    => dsp0_d_i(3)
   ,  D5    => dsp0_d_i(4)
   ,  D6    => dsp0_d_i(5)
   ,  D7    => dsp0_d_i(6)
   ,  D8    => dsp0_d_i(7)
   ,  D9    => dsp0_d_i(8)
   ,  D10   => dsp0_d_i(9)
   ,  D11   => dsp0_d_i(10)
   ,  D12   => dsp0_d_i(11)
   ,  D13   => dsp0_d_i(12)
   ,  D14   => dsp0_d_i(13)
   ,  D15   => dsp0_d_i(14)
   ,  D16   => dsp0_d_i(15)
   ,  D17   => dsp0_d_i(16)
   ,  D18   => dsp0_d_i(17)
   ,  OVF   => dsp0_ovf_o
   ,  R     => dsp0_rst_i
   ,  RZ    => dsp0_rstz_i
   ,  WE    => dsp0_we_i
   ,  Z1    => dsp0_z_o(0)
   ,  Z2    => dsp0_z_o(1)
   ,  Z3    => dsp0_z_o(2)
   ,  Z4    => dsp0_z_o(3)
   ,  Z5    => dsp0_z_o(4)
   ,  Z6    => dsp0_z_o(5)
   ,  Z7    => dsp0_z_o(6)
   ,  Z8    => dsp0_z_o(7)
   ,  Z9    => dsp0_z_o(8)
   ,  Z10   => dsp0_z_o(9)
   ,  Z11   => dsp0_z_o(10)
   ,  Z12   => dsp0_z_o(11)
   ,  Z13   => dsp0_z_o(12)
   ,  Z14   => dsp0_z_o(13)
   ,  Z15   => dsp0_z_o(14)
   ,  Z16   => dsp0_z_o(15)
   ,  Z17   => dsp0_z_o(16)
   ,  Z18   => dsp0_z_o(17)
   ,  Z19   => dsp0_z_o(18)
   ,  Z20   => dsp0_z_o(19)
   ,  Z21   => dsp0_z_o(20)
   ,  Z22   => dsp0_z_o(21)
   ,  Z23   => dsp0_z_o(22)
   ,  Z24   => dsp0_z_o(23)
   ,  Z25   => dsp0_z_o(24)
   ,  Z26   => dsp0_z_o(25)
   ,  Z27   => dsp0_z_o(26)
   ,  Z28   => dsp0_z_o(27)
   ,  Z29   => dsp0_z_o(28)
   ,  Z30   => dsp0_z_o(29)
   ,  Z31   => dsp0_z_o(30)
   ,  Z32   => dsp0_z_o(31)
   ,  Z33   => dsp0_z_o(32)
   ,  Z34   => dsp0_z_o(33)
   ,  Z35   => dsp0_z_o(34)
   ,  Z36   => dsp0_z_o(35)
   ,  Z37   => dsp0_z_o(36)
   ,  Z38   => dsp0_z_o(37)
   ,  Z39   => dsp0_z_o(38)
   ,  Z40   => dsp0_z_o(39)
   ,  Z41   => dsp0_z_o(40)
   ,  Z42   => dsp0_z_o(41)
   ,  Z43   => dsp0_z_o(42)
   ,  Z44   => dsp0_z_o(43)
   ,  Z45   => dsp0_z_o(44)
   ,  Z46   => dsp0_z_o(45)
   ,  Z47   => dsp0_z_o(46)
   ,  Z48   => dsp0_z_o(47)
   ,  Z49   => dsp0_z_o(48)
   ,  Z50   => dsp0_z_o(49)
   ,  Z51   => dsp0_z_o(50)
   ,  Z52   => dsp0_z_o(51)
   ,  Z53   => dsp0_z_o(52)
   ,  Z54   => dsp0_z_o(53)
   ,  Z55   => dsp0_z_o(54)
   ,  Z56   => dsp0_z_o(55)
);
--#}}}#

-- instance dsp1#{{{#
dsp_1 : NX_DSP_L_BOX
generic map (
    col    => col
  , row    => row
  , cfg0_i => cfg0_i
  , cfg1_i => cfg1_i
)
port map (
      A1    => dsp1_a_i(0)
   ,  A2    => dsp1_a_i(1)
   ,  A3    => dsp1_a_i(2)
   ,  A4    => dsp1_a_i(3)
   ,  A5    => dsp1_a_i(4)
   ,  A6    => dsp1_a_i(5)
   ,  A7    => dsp1_a_i(6)
   ,  A8    => dsp1_a_i(7)
   ,  A9    => dsp1_a_i(8)
   ,  A10   => dsp1_a_i(9)
   ,  A11   => dsp1_a_i(10)
   ,  A12   => dsp1_a_i(11)
   ,  A13   => dsp1_a_i(12)
   ,  A14   => dsp1_a_i(13)
   ,  A15   => dsp1_a_i(14)
   ,  A16   => dsp1_a_i(15)
   ,  A17   => dsp1_a_i(16)
   ,  A18   => dsp1_a_i(17)
   ,  A19   => dsp1_a_i(18)
   ,  A20   => dsp1_a_i(19)
   ,  A21   => dsp1_a_i(20)
   ,  A22   => dsp1_a_i(21)
   ,  A23   => dsp1_a_i(22)
   ,  A24   => dsp1_a_i(23)
   ,  B1    => dsp1_b_i(0)
   ,  B2    => dsp1_b_i(1)
   ,  B3    => dsp1_b_i(2)
   ,  B4    => dsp1_b_i(3)
   ,  B5    => dsp1_b_i(4)
   ,  B6    => dsp1_b_i(5)
   ,  B7    => dsp1_b_i(6)
   ,  B8    => dsp1_b_i(7)
   ,  B9    => dsp1_b_i(8)
   ,  B10   => dsp1_b_i(9)
   ,  B11   => dsp1_b_i(10)
   ,  B12   => dsp1_b_i(11)
   ,  B13   => dsp1_b_i(12)
   ,  B14   => dsp1_b_i(13)
   ,  B15   => dsp1_b_i(14)
   ,  B16   => dsp1_b_i(15)
   ,  B17   => dsp1_b_i(16)
   ,  B18   => dsp1_b_i(17)
   ,  C1    => dsp1_c_i(0)
   ,  C2    => dsp1_c_i(1)
   ,  C3    => dsp1_c_i(2)
   ,  C4    => dsp1_c_i(3)
   ,  C5    => dsp1_c_i(4)
   ,  C6    => dsp1_c_i(5)
   ,  C7    => dsp1_c_i(6)
   ,  C8    => dsp1_c_i(7)
   ,  C9    => dsp1_c_i(8)
   ,  C10   => dsp1_c_i(9)
   ,  C11   => dsp1_c_i(10)
   ,  C12   => dsp1_c_i(11)
   ,  C13   => dsp1_c_i(12)
   ,  C14   => dsp1_c_i(13)
   ,  C15   => dsp1_c_i(14)
   ,  C16   => dsp1_c_i(15)
   ,  C17   => dsp1_c_i(16)
   ,  C18   => dsp1_c_i(17)
   ,  C19   => dsp1_c_i(18)
   ,  C20   => dsp1_c_i(19)
   ,  C21   => dsp1_c_i(20)
   ,  C22   => dsp1_c_i(21)
   ,  C23   => dsp1_c_i(22)
   ,  C24   => dsp1_c_i(23)
   ,  C25   => dsp1_c_i(24)
   ,  C26   => dsp1_c_i(25)
   ,  C27   => dsp1_c_i(26)
   ,  C28   => dsp1_c_i(27)
   ,  C29   => dsp1_c_i(28)
   ,  C30   => dsp1_c_i(29)
   ,  C31   => dsp1_c_i(30)
   ,  C32   => dsp1_c_i(31)
   ,  C33   => dsp1_c_i(32)
   ,  C34   => dsp1_c_i(33)
   ,  C35   => dsp1_c_i(34)
   ,  C36   => dsp1_c_i(35)
   ,  CAI1  => dsp_ca_i(0)
   ,  CAI2  => dsp_ca_i(1)
   ,  CAI3  => dsp_ca_i(2)
   ,  CAI4  => dsp_ca_i(3)
   ,  CAI5  => dsp_ca_i(4)
   ,  CAI6  => dsp_ca_i(5)
   ,  CAI7  => dsp_ca_i(6)
   ,  CAI8  => dsp_ca_i(7)
   ,  CAI9  => dsp_ca_i(8)
   ,  CAI10 => dsp_ca_i(9)
   ,  CAI11 => dsp_ca_i(10)
   ,  CAI12 => dsp_ca_i(11)
   ,  CAI13 => dsp_ca_i(12)
   ,  CAI14 => dsp_ca_i(13)
   ,  CAI15 => dsp_ca_i(14)
   ,  CAI16 => dsp_ca_i(15)
   ,  CAI17 => dsp_ca_i(16)
   ,  CAI18 => dsp_ca_i(17)
   ,  CAI19 => dsp_ca_i(18)
   ,  CAI20 => dsp_ca_i(19)
   ,  CAI21 => dsp_ca_i(20)
   ,  CAI22 => dsp_ca_i(21)
   ,  CAI23 => dsp_ca_i(22)
   ,  CAI24 => dsp_ca_i(23)
   ,  CAO1  => c_a_int(0)
   ,  CAO2  => c_a_int(1)
   ,  CAO3  => c_a_int(2)
   ,  CAO4  => c_a_int(3)
   ,  CAO5  => c_a_int(4)
   ,  CAO6  => c_a_int(5)
   ,  CAO7  => c_a_int(6)
   ,  CAO8  => c_a_int(7)
   ,  CAO9  => c_a_int(8)
   ,  CAO10 => c_a_int(9)
   ,  CAO11 => c_a_int(10)
   ,  CAO12 => c_a_int(11)
   ,  CAO13 => c_a_int(12)
   ,  CAO14 => c_a_int(13)
   ,  CAO15 => c_a_int(14)
   ,  CAO16 => c_a_int(15)
   ,  CAO17 => c_a_int(16)
   ,  CAO18 => c_a_int(17)
   ,  CAO19 => c_a_int(18)
   ,  CAO20 => c_a_int(19)
   ,  CAO21 => c_a_int(20)
   ,  CAO22 => c_a_int(21)
   ,  CAO23 => c_a_int(22)
   ,  CAO24 => c_a_int(23)
   ,  CBI1  => dsp_cb_i(0)
   ,  CBI2  => dsp_cb_i(1)
   ,  CBI3  => dsp_cb_i(2)
   ,  CBI4  => dsp_cb_i(3)
   ,  CBI5  => dsp_cb_i(4)
   ,  CBI6  => dsp_cb_i(5)
   ,  CBI7  => dsp_cb_i(6)
   ,  CBI8  => dsp_cb_i(7)
   ,  CBI9  => dsp_cb_i(8)
   ,  CBI10 => dsp_cb_i(9)
   ,  CBI11 => dsp_cb_i(10)
   ,  CBI12 => dsp_cb_i(11)
   ,  CBI13 => dsp_cb_i(12)
   ,  CBI14 => dsp_cb_i(13)
   ,  CBI15 => dsp_cb_i(14)
   ,  CBI16 => dsp_cb_i(15)
   ,  CBI17 => dsp_cb_i(16)
   ,  CBI18 => dsp_cb_i(17)
   ,  CBO1  => c_b_int(0)
   ,  CBO2  => c_b_int(1)
   ,  CBO3  => c_b_int(2)
   ,  CBO4  => c_b_int(3)
   ,  CBO5  => c_b_int(4)
   ,  CBO6  => c_b_int(5)
   ,  CBO7  => c_b_int(6)
   ,  CBO8  => c_b_int(7)
   ,  CBO9  => c_b_int(8)
   ,  CBO10 => c_b_int(9)
   ,  CBO11 => c_b_int(10)
   ,  CBO12 => c_b_int(11)
   ,  CBO13 => c_b_int(12)
   ,  CBO14 => c_b_int(13)
   ,  CBO15 => c_b_int(14)
   ,  CBO16 => c_b_int(15)
   ,  CBO17 => c_b_int(16)
   ,  CBO18 => c_b_int(17)
   ,  CCI   => c_cy_int
   ,  CCO   => dsp_ccy_o
   ,  CI    => dsp1_cy_i
   ,  CK    => dsp1_clk_i
   ,  CO    => dsp1_cy_o
   ,  CO37  => dsp1_cy36_o
   ,  CO57  => dsp1_cy56_o
   ,  CZI1  => dsp_cz_i(0)
   ,  CZI2  => dsp_cz_i(1)
   ,  CZI3  => dsp_cz_i(2)
   ,  CZI4  => dsp_cz_i(3)
   ,  CZI5  => dsp_cz_i(4)
   ,  CZI6  => dsp_cz_i(5)
   ,  CZI7  => dsp_cz_i(6)
   ,  CZI8  => dsp_cz_i(7)
   ,  CZI9  => dsp_cz_i(8)
   ,  CZI10 => dsp_cz_i(9)
   ,  CZI11 => dsp_cz_i(10)
   ,  CZI12 => dsp_cz_i(11)
   ,  CZI13 => dsp_cz_i(12)
   ,  CZI14 => dsp_cz_i(13)
   ,  CZI15 => dsp_cz_i(14)
   ,  CZI16 => dsp_cz_i(15)
   ,  CZI17 => dsp_cz_i(16)
   ,  CZI18 => dsp_cz_i(17)
   ,  CZI19 => dsp_cz_i(18)
   ,  CZI20 => dsp_cz_i(19)
   ,  CZI21 => dsp_cz_i(20)
   ,  CZI22 => dsp_cz_i(21)
   ,  CZI23 => dsp_cz_i(22)
   ,  CZI24 => dsp_cz_i(23)
   ,  CZI25 => dsp_cz_i(24)
   ,  CZI26 => dsp_cz_i(25)
   ,  CZI27 => dsp_cz_i(26)
   ,  CZI28 => dsp_cz_i(27)
   ,  CZI29 => dsp_cz_i(28)
   ,  CZI30 => dsp_cz_i(29)
   ,  CZI31 => dsp_cz_i(30)
   ,  CZI32 => dsp_cz_i(31)
   ,  CZI33 => dsp_cz_i(32)
   ,  CZI34 => dsp_cz_i(33)
   ,  CZI35 => dsp_cz_i(34)
   ,  CZI36 => dsp_cz_i(35)
   ,  CZI37 => dsp_cz_i(36)
   ,  CZI38 => dsp_cz_i(37)
   ,  CZI39 => dsp_cz_i(38)
   ,  CZI40 => dsp_cz_i(39)
   ,  CZI41 => dsp_cz_i(40)
   ,  CZI42 => dsp_cz_i(41)
   ,  CZI43 => dsp_cz_i(42)
   ,  CZI44 => dsp_cz_i(43)
   ,  CZI45 => dsp_cz_i(44)
   ,  CZI46 => dsp_cz_i(45)
   ,  CZI47 => dsp_cz_i(46)
   ,  CZI48 => dsp_cz_i(47)
   ,  CZI49 => dsp_cz_i(48)
   ,  CZI50 => dsp_cz_i(49)
   ,  CZI51 => dsp_cz_i(50)
   ,  CZI52 => dsp_cz_i(51)
   ,  CZI53 => dsp_cz_i(52)
   ,  CZI54 => dsp_cz_i(53)
   ,  CZI55 => dsp_cz_i(54)
   ,  CZI56 => dsp_cz_i(55)
   ,  CZO1  => c_z_int(0)
   ,  CZO2  => c_z_int(1)
   ,  CZO3  => c_z_int(2)
   ,  CZO4  => c_z_int(3)
   ,  CZO5  => c_z_int(4)
   ,  CZO6  => c_z_int(5)
   ,  CZO7  => c_z_int(6)
   ,  CZO8  => c_z_int(7)
   ,  CZO9  => c_z_int(8)
   ,  CZO10 => c_z_int(9)
   ,  CZO11 => c_z_int(10)
   ,  CZO12 => c_z_int(11)
   ,  CZO13 => c_z_int(12)
   ,  CZO14 => c_z_int(13)
   ,  CZO15 => c_z_int(14)
   ,  CZO16 => c_z_int(15)
   ,  CZO17 => c_z_int(16)
   ,  CZO18 => c_z_int(17)
   ,  CZO19 => c_z_int(18)
   ,  CZO20 => c_z_int(19)
   ,  CZO21 => c_z_int(20)
   ,  CZO22 => c_z_int(21)
   ,  CZO23 => c_z_int(22)
   ,  CZO24 => c_z_int(23)
   ,  CZO25 => c_z_int(24)
   ,  CZO26 => c_z_int(25)
   ,  CZO27 => c_z_int(26)
   ,  CZO28 => c_z_int(27)
   ,  CZO29 => c_z_int(28)
   ,  CZO30 => c_z_int(29)
   ,  CZO31 => c_z_int(30)
   ,  CZO32 => c_z_int(31)
   ,  CZO33 => c_z_int(32)
   ,  CZO34 => c_z_int(33)
   ,  CZO35 => c_z_int(34)
   ,  CZO36 => c_z_int(35)
   ,  CZO37 => c_z_int(36)
   ,  CZO38 => c_z_int(37)
   ,  CZO39 => c_z_int(38)
   ,  CZO40 => c_z_int(39)
   ,  CZO41 => c_z_int(40)
   ,  CZO42 => c_z_int(41)
   ,  CZO43 => c_z_int(42)
   ,  CZO44 => c_z_int(43)
   ,  CZO45 => c_z_int(44)
   ,  CZO46 => c_z_int(45)
   ,  CZO47 => c_z_int(46)
   ,  CZO48 => c_z_int(47)
   ,  CZO49 => c_z_int(48)
   ,  CZO50 => c_z_int(49)
   ,  CZO51 => c_z_int(50)
   ,  CZO52 => c_z_int(51)
   ,  CZO53 => c_z_int(52)
   ,  CZO54 => c_z_int(53)
   ,  CZO55 => c_z_int(54)
   ,  CZO56 => c_z_int(55)
   ,  D1    => dsp1_d_i(0)
   ,  D2    => dsp1_d_i(1)
   ,  D3    => dsp1_d_i(2)
   ,  D4    => dsp1_d_i(3)
   ,  D5    => dsp1_d_i(4)
   ,  D6    => dsp1_d_i(5)
   ,  D7    => dsp1_d_i(6)
   ,  D8    => dsp1_d_i(7)
   ,  D9    => dsp1_d_i(8)
   ,  D10   => dsp1_d_i(9)
   ,  D11   => dsp1_d_i(10)
   ,  D12   => dsp1_d_i(11)
   ,  D13   => dsp1_d_i(12)
   ,  D14   => dsp1_d_i(13)
   ,  D15   => dsp1_d_i(14)
   ,  D16   => dsp1_d_i(15)
   ,  D17   => dsp1_d_i(16)
   ,  D18   => dsp1_d_i(17)
   ,  OVF   => dsp1_ovf_o
   ,  R     => dsp1_rst_i
   ,  RZ    => dsp1_rstz_i
   ,  WE    => dsp1_we_i
   ,  Z1    => dsp1_z_o(0)
   ,  Z2    => dsp1_z_o(1)
   ,  Z3    => dsp1_z_o(2)
   ,  Z4    => dsp1_z_o(3)
   ,  Z5    => dsp1_z_o(4)
   ,  Z6    => dsp1_z_o(5)
   ,  Z7    => dsp1_z_o(6)
   ,  Z8    => dsp1_z_o(7)
   ,  Z9    => dsp1_z_o(8)
   ,  Z10   => dsp1_z_o(9)
   ,  Z11   => dsp1_z_o(10)
   ,  Z12   => dsp1_z_o(11)
   ,  Z13   => dsp1_z_o(12)
   ,  Z14   => dsp1_z_o(13)
   ,  Z15   => dsp1_z_o(14)
   ,  Z16   => dsp1_z_o(15)
   ,  Z17   => dsp1_z_o(16)
   ,  Z18   => dsp1_z_o(17)
   ,  Z19   => dsp1_z_o(18)
   ,  Z20   => dsp1_z_o(19)
   ,  Z21   => dsp1_z_o(20)
   ,  Z22   => dsp1_z_o(21)
   ,  Z23   => dsp1_z_o(22)
   ,  Z24   => dsp1_z_o(23)
   ,  Z25   => dsp1_z_o(24)
   ,  Z26   => dsp1_z_o(25)
   ,  Z27   => dsp1_z_o(26)
   ,  Z28   => dsp1_z_o(27)
   ,  Z29   => dsp1_z_o(28)
   ,  Z30   => dsp1_z_o(29)
   ,  Z31   => dsp1_z_o(30)
   ,  Z32   => dsp1_z_o(31)
   ,  Z33   => dsp1_z_o(32)
   ,  Z34   => dsp1_z_o(33)
   ,  Z35   => dsp1_z_o(34)
   ,  Z36   => dsp1_z_o(35)
   ,  Z37   => dsp1_z_o(36)
   ,  Z38   => dsp1_z_o(37)
   ,  Z39   => dsp1_z_o(38)
   ,  Z40   => dsp1_z_o(39)
   ,  Z41   => dsp1_z_o(40)
   ,  Z42   => dsp1_z_o(41)
   ,  Z43   => dsp1_z_o(42)
   ,  Z44   => dsp1_z_o(43)
   ,  Z45   => dsp1_z_o(44)
   ,  Z46   => dsp1_z_o(45)
   ,  Z47   => dsp1_z_o(46)
   ,  Z48   => dsp1_z_o(47)
   ,  Z49   => dsp1_z_o(48)
   ,  Z50   => dsp1_z_o(49)
   ,  Z51   => dsp1_z_o(50)
   ,  Z52   => dsp1_z_o(51)
   ,  Z53   => dsp1_z_o(52)
   ,  Z54   => dsp1_z_o(53)
   ,  Z55   => dsp1_z_o(54)
   ,  Z56   => dsp1_z_o(55)
);
--#}}}#

-- instance ram0#{{{#
ram_0 : NX_RAM_L_BOX
generic map (
    col    => col
  , row    => row
  , cfg0_i => cfg0_i
  , cfg1_i => cfg1_i
)
port map (
    ACK   => dpram_clkmem0_i
  , ACKC  => dpram_clkmemclone0_i
  , ACKD  => dpram_clkmem90_0_i
  , ACKR  => dpram_clkreg0_i
  , BCK   => dpram_clkmem1_i
  , BCKC  => dpram_clkmemclone1_i
  , BCKD  => dpram_clkmem90_1_i
  , BCKR  => dpram_clkreg1_i

  , AI1   => dpram_din0_i(0)
  , AI2   => dpram_din0_i(1)
  , AI3   => dpram_din0_i(2)
  , AI4   => dpram_din0_i(3)
  , AI5   => dpram_din0_i(4)
  , AI6   => dpram_din0_i(5)
  , AI7   => dpram_din0_i(6)
  , AI8   => dpram_din0_i(7)
  , AI9   => dpram_din0_i(8)
  , AI10  => dpram_din0_i(9)
  , AI11  => dpram_din0_i(10)
  , AI12  => dpram_din0_i(11)
  , AI13  => dpram_din0_i(12)
  , AI14  => dpram_din0_i(13)
  , AI15  => dpram_din0_i(14)
  , AI16  => dpram_din0_i(15)
  , AI17  => dpram_din0_i(16)
  , AI18  => dpram_din0_i(17)
  , AI19  => dpram_din0_i(18)
  , AI20  => dpram_din0_i(19)
  , AI21  => dpram_din0_i(20)
  , AI22  => dpram_din0_i(21)
  , AI23  => dpram_din0_i(22)
  , AI24  => dpram_din0_i(23)

  , BI1   => dpram_din1_i(0)
  , BI2   => dpram_din1_i(1)
  , BI3   => dpram_din1_i(2)
  , BI4   => dpram_din1_i(3)
  , BI5   => dpram_din1_i(4)
  , BI6   => dpram_din1_i(5)
  , BI7   => dpram_din1_i(6)
  , BI8   => dpram_din1_i(7)
  , BI9   => dpram_din1_i(8)
  , BI10  => dpram_din1_i(9)
  , BI11  => dpram_din1_i(10)
  , BI12  => dpram_din1_i(11)
  , BI13  => dpram_din1_i(12)
  , BI14  => dpram_din1_i(13)
  , BI15  => dpram_din1_i(14)
  , BI16  => dpram_din1_i(15)
  , BI17  => dpram_din1_i(16)
  , BI18  => dpram_din1_i(17)
  , BI19  => dpram_din1_i(18)
  , BI20  => dpram_din1_i(19)
  , BI21  => dpram_din1_i(20)
  , BI22  => dpram_din1_i(21)
  , BI23  => dpram_din1_i(22)
  , BI24  => dpram_din1_i(23)

  , ACOR => dpram_ecc_corrected0_o
  , AERR => dpram_ecc_uncorrected0_o
  , BCOR => dpram_ecc_corrected1_o
  , BERR => dpram_ecc_uncorrected1_o

  , AO1  => dpram_dout0_o(0)
  , AO2  => dpram_dout0_o(1)
  , AO3  => dpram_dout0_o(2)
  , AO4  => dpram_dout0_o(3)
  , AO5  => dpram_dout0_o(4)
  , AO6  => dpram_dout0_o(5)
  , AO7  => dpram_dout0_o(6)
  , AO8  => dpram_dout0_o(7)
  , AO9  => dpram_dout0_o(8)
  , AO10 => dpram_dout0_o(9)
  , AO11 => dpram_dout0_o(10)
  , AO12 => dpram_dout0_o(11)
  , AO13 => dpram_dout0_o(12)
  , AO14 => dpram_dout0_o(13)
  , AO15 => dpram_dout0_o(14)
  , AO16 => dpram_dout0_o(15)
  , AO17 => dpram_dout0_o(16)
  , AO18 => dpram_dout0_o(17)
  , AO19 => dpram_dout0_o(18)
  , AO20 => dpram_dout0_o(19)
  , AO21 => dpram_dout0_o(20)
  , AO22 => dpram_dout0_o(21)
  , AO23 => dpram_dout0_o(22)
  , AO24 => dpram_dout0_o(23)

  , BO1  => dpram_dout1_o(0)
  , BO2  => dpram_dout1_o(1)
  , BO3  => dpram_dout1_o(2)
  , BO4  => dpram_dout1_o(3)
  , BO5  => dpram_dout1_o(4)
  , BO6  => dpram_dout1_o(5)
  , BO7  => dpram_dout1_o(6)
  , BO8  => dpram_dout1_o(7)
  , BO9  => dpram_dout1_o(8)
  , BO10 => dpram_dout1_o(9)
  , BO11 => dpram_dout1_o(10)
  , BO12 => dpram_dout1_o(11)
  , BO13 => dpram_dout1_o(12)
  , BO14 => dpram_dout1_o(13)
  , BO15 => dpram_dout1_o(14)
  , BO16 => dpram_dout1_o(15)
  , BO17 => dpram_dout1_o(16)
  , BO18 => dpram_dout1_o(17)
  , BO19 => dpram_dout1_o(18)
  , BO20 => dpram_dout1_o(19)
  , BO21 => dpram_dout1_o(20)
  , BO22 => dpram_dout1_o(21)
  , BO23 => dpram_dout1_o(22)
  , BO24 => dpram_dout1_o(23)

  , AA1  => dpram_addr0_i(0)
  , AA2  => dpram_addr0_i(1)
  , AA3  => dpram_addr0_i(2)
  , AA4  => dpram_addr0_i(3)
  , AA5  => dpram_addr0_i(4)
  , AA6  => dpram_addr0_i(5)
  , AA7  => dpram_addr0_i(6)
  , AA8  => dpram_addr0_i(7)
  , AA9  => dpram_addr0_i(8)
  , AA10 => dpram_addr0_i(9)
  , AA11 => dpram_addr0_i(10)
  , AA12 => dpram_addr0_i(11)
  , AA13 => dpram_addr0_i(12)
  , AA14 => dpram_addr0_i(13)
  , AA15 => dpram_addr0_i(14)
  , AA16 => dpram_addr0_i(15)

  , ACS  => dpram_cs0_i
  , AWE  => dpram_we0_i
  , AR   => dpram_rst0_i

  , BA1  => dpram_addr1_i(0)
  , BA2  => dpram_addr1_i(1)
  , BA3  => dpram_addr1_i(2)
  , BA4  => dpram_addr1_i(3)
  , BA5  => dpram_addr1_i(4)
  , BA6  => dpram_addr1_i(5)
  , BA7  => dpram_addr1_i(6)
  , BA8  => dpram_addr1_i(7)
  , BA9  => dpram_addr1_i(8)
  , BA10 => dpram_addr1_i(9)
  , BA11 => dpram_addr1_i(10)
  , BA12 => dpram_addr1_i(11)
  , BA13 => dpram_addr1_i(12)
  , BA14 => dpram_addr1_i(13)
  , BA15 => dpram_addr1_i(14)
  , BA16 => dpram_addr1_i(15)

  , BCS  => dpram_cs1_i
  , BWE  => dpram_we1_i
  , BR   => dpram_rst1_i
);
--#}}}#

end NX_RTL;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_L_BOX definition
-- =================================================================================================

-- NX_DSP_L_BOX#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_DSP_L_BOX is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end NX_DSP_L_BOX;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RAM_L_BOX definition
-- =================================================================================================

-- NX_RAM_L_BOX #{{{#
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_RAM_L_BOX is
generic (
    col    : integer := 2;
    row    : integer := 4;
    cfg0_i : bit_vector(95 downto 0) := (others => '0');
    cfg1_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    ACK   : in  std_logic;
    ACKC  : in  std_logic;
    ACKD  : in  std_logic;
    ACKR  : in  std_logic;
    BCK   : in  std_logic;
    BCKC  : in  std_logic;
    BCKD  : in  std_logic;
    BCKR  : in  std_logic;

    AI1   : in  std_logic;
    AI2   : in  std_logic;
    AI3   : in  std_logic;
    AI4   : in  std_logic;
    AI5   : in  std_logic;
    AI6   : in  std_logic;
    AI7   : in  std_logic;
    AI8   : in  std_logic;
    AI9   : in  std_logic;
    AI10  : in  std_logic;
    AI11  : in  std_logic;
    AI12  : in  std_logic;
    AI13  : in  std_logic;
    AI14  : in  std_logic;
    AI15  : in  std_logic;
    AI16  : in  std_logic;

    AI17  : in  std_logic;
    AI18  : in  std_logic;
    AI19  : in  std_logic;
    AI20  : in  std_logic;
    AI21  : in  std_logic;
    AI22  : in  std_logic;
    AI23  : in  std_logic;
    AI24  : in  std_logic;

    BI1   : in  std_logic;
    BI2   : in  std_logic;
    BI3   : in  std_logic;
    BI4   : in  std_logic;
    BI5   : in  std_logic;
    BI6   : in  std_logic;
    BI7   : in  std_logic;
    BI8   : in  std_logic;
    BI9   : in  std_logic;
    BI10  : in  std_logic;
    BI11  : in  std_logic;
    BI12  : in  std_logic;
    BI13  : in  std_logic;
    BI14  : in  std_logic;
    BI15  : in  std_logic;
    BI16  : in  std_logic;

    BI17  : in  std_logic;
    BI18  : in  std_logic;
    BI19  : in  std_logic;
    BI20  : in  std_logic;
    BI21  : in  std_logic;
    BI22  : in  std_logic;
    BI23  : in  std_logic;
    BI24  : in  std_logic;

    ACOR  : out std_logic;
    AERR  : out std_logic;
    BCOR  : out std_logic;
    BERR  : out std_logic;

    AO1   : out std_logic;
    AO2   : out std_logic;
    AO3   : out std_logic;
    AO4   : out std_logic;
    AO5   : out std_logic;
    AO6   : out std_logic;
    AO7   : out std_logic;
    AO8   : out std_logic;
    AO9   : out std_logic;
    AO10  : out std_logic;
    AO11  : out std_logic;
    AO12  : out std_logic;
    AO13  : out std_logic;
    AO14  : out std_logic;
    AO15  : out std_logic;
    AO16  : out std_logic;

    AO17  : out std_logic;
    AO18  : out std_logic;
    AO19  : out std_logic;
    AO20  : out std_logic;
    AO21  : out std_logic;
    AO22  : out std_logic;
    AO23  : out std_logic;
    AO24  : out std_logic;

    BO1   : out std_logic;
    BO2   : out std_logic;
    BO3   : out std_logic;
    BO4   : out std_logic;
    BO5   : out std_logic;
    BO6   : out std_logic;
    BO7   : out std_logic;
    BO8   : out std_logic;
    BO9   : out std_logic;
    BO10  : out std_logic;
    BO11  : out std_logic;
    BO12  : out std_logic;
    BO13  : out std_logic;
    BO14  : out std_logic;
    BO15  : out std_logic;
    BO16  : out std_logic;

    BO17  : out std_logic;
    BO18  : out std_logic;
    BO19  : out std_logic;
    BO20  : out std_logic;
    BO21  : out std_logic;
    BO22  : out std_logic;
    BO23  : out std_logic;
    BO24  : out std_logic;

    AA1   : in  std_logic;
    AA2   : in  std_logic;
    AA3   : in  std_logic;
    AA4   : in  std_logic;
    AA5   : in  std_logic;
    AA6   : in  std_logic;

    AA7   : in  std_logic;
    AA8   : in  std_logic;
    AA9   : in  std_logic;
    AA10  : in  std_logic;
    AA11  : in  std_logic;
    AA12  : in  std_logic;
    AA13  : in  std_logic;
    AA14  : in  std_logic;
    AA15  : in  std_logic;
    AA16  : in  std_logic;

    ACS   : in  std_logic;
    AWE   : in  std_logic;
    AR    : in  std_logic;

    BA1   : in  std_logic;
    BA2   : in  std_logic;
    BA3   : in  std_logic;
    BA4   : in  std_logic;
    BA5   : in  std_logic;
    BA6   : in  std_logic;

    BA7   : in  std_logic;
    BA8   : in  std_logic;
    BA9   : in  std_logic;
    BA10  : in  std_logic;
    BA11  : in  std_logic;
    BA12  : in  std_logic;
    BA13  : in  std_logic;
    BA14  : in  std_logic;
    BA15  : in  std_logic;
    BA16  : in  std_logic;

    BCS   : in  std_logic;
    BWE   : in  std_logic;
    BR    : in  std_logic
);
end NX_RAM_L_BOX;
--#}}}}
-- =================================================================================================
--   NX_DSP_L definition                                                                2018/11/30
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DSP_L is
generic (
    std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";   -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";    -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";          -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                 -- ALU
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end NX_DSP_L;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_L_WRAP definition                                                           2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity NX_DSP_L_WRAP is
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A    : in  std_logic_vector(23 downto 0);
    B    : in  std_logic_vector(17 downto 0);
    C    : in  std_logic_vector(35 downto 0);

    CAI  : in  std_logic_vector(23 downto 0);
    CAO  : out std_logic_vector(23 downto 0);
    CBI  : in  std_logic_vector(17 downto 0);
    CBO  : out std_logic_vector(17 downto 0);

    CCI  : in  std_logic;
    CCO  : out std_logic;
    CI   : in  std_logic;
    CK   : in  std_logic;
    CO   : out std_logic;
    CO37 : out std_logic;
    CO57 : out std_logic;

    CZI  : in  std_logic_vector(55 downto 0);
    CZO  : out std_logic_vector(55 downto 0);

    D    : in  std_logic_vector(17 downto 0);

    OVF  : out std_logic;
    R    : in  std_logic;
    RZ   : in  std_logic;
    WE   : in  std_logic;

    Z    : out std_logic_vector(55 downto 0)
);
end NX_DSP_L_WRAP;

-- architecture NX_ARCH of NX_DSP_L_WRAP#{{{#
architecture NX_ARCH of NX_DSP_L_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_ARCH: architecture is "WRAPPER";

component NX_DSP_L
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";      -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";       -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";             -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                    -- ALU
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end component;

begin

dsp: NX_DSP_L generic map (
    std_mode    => std_mode,
    raw_config0 => raw_config0,
    raw_config1 => raw_config1,
    raw_config2 => raw_config2,
    raw_config3 => raw_config3)
port map (
    A1    => A(0),
    A2    => A(1),
    A3    => A(2),
    A4    => A(3),
    A5    => A(4),
    A6    => A(5),
    A7    => A(6),
    A8    => A(7),
    A9    => A(8),
    A10   => A(9),
    A11   => A(10),
    A12   => A(11),
    A13   => A(12),
    A14   => A(13),
    A15   => A(14),
    A16   => A(15),
    A17   => A(16),
    A18   => A(17),
    A19   => A(18),
    A20   => A(19),
    A21   => A(20),
    A22   => A(21),
    A23   => A(22),
    A24   => A(23),

    B1    => B(0),
    B2    => B(1),
    B3    => B(2),
    B4    => B(3),
    B5    => B(4),
    B6    => B(5),
    B7    => B(6),
    B8    => B(7),
    B9    => B(8),
    B10   => B(9),
    B11   => B(10),
    B12   => B(11),
    B13   => B(12),
    B14   => B(13),
    B15   => B(14),
    B16   => B(15),
    B17   => B(16),
    B18   => B(17),

    C1    => C(0),
    C2    => C(1),
    C3    => C(2),
    C4    => C(3),
    C5    => C(4),
    C6    => C(5),
    C7    => C(6),
    C8    => C(7),
    C9    => C(8),
    C10   => C(9),
    C11   => C(10),
    C12   => C(11),
    C13   => C(12),
    C14   => C(13),
    C15   => C(14),
    C16   => C(15),
    C17   => C(16),
    C18   => C(17),
    C19   => C(18),
    C20   => C(19),
    C21   => C(20),
    C22   => C(21),
    C23   => C(22),
    C24   => C(23),
    C25   => C(24),
    C26   => C(25),
    C27   => C(26),
    C28   => C(27),
    C29   => C(28),
    C30   => C(29),
    C31   => C(30),
    C32   => C(31),
    C33   => C(32),
    C34   => C(33),
    C35   => C(34),
    C36   => C(35),

    CAI1  => CAI(0),
    CAI2  => CAI(1),
    CAI3  => CAI(2),
    CAI4  => CAI(3),
    CAI5  => CAI(4),
    CAI6  => CAI(5),
    CAI7  => CAI(6),
    CAI8  => CAI(7),
    CAI9  => CAI(8),
    CAI10 => CAI(9),
    CAI11 => CAI(10),
    CAI12 => CAI(11),
    CAI13 => CAI(12),
    CAI14 => CAI(13),
    CAI15 => CAI(14),
    CAI16 => CAI(15),
    CAI17 => CAI(16),
    CAI18 => CAI(17),
    CAI19 => CAI(18),
    CAI20 => CAI(19),
    CAI21 => CAI(20),
    CAI22 => CAI(21),
    CAI23 => CAI(22),
    CAI24 => CAI(23),

    CAO1  => CAO(0),
    CAO2  => CAO(1),
    CAO3  => CAO(2),
    CAO4  => CAO(3),
    CAO5  => CAO(4),
    CAO6  => CAO(5),
    CAO7  => CAO(6),
    CAO8  => CAO(7),
    CAO9  => CAO(8),
    CAO10 => CAO(9),
    CAO11 => CAO(10),
    CAO12 => CAO(11),
    CAO13 => CAO(12),
    CAO14 => CAO(13),
    CAO15 => CAO(14),
    CAO16 => CAO(15),
    CAO17 => CAO(16),
    CAO18 => CAO(17),
    CAO19 => CAO(18),
    CAO20 => CAO(19),
    CAO21 => CAO(20),
    CAO22 => CAO(21),
    CAO23 => CAO(22),
    CAO24 => CAO(23),

    CBI1  => CBI(0),
    CBI2  => CBI(1),
    CBI3  => CBI(2),
    CBI4  => CBI(3),
    CBI5  => CBI(4),
    CBI6  => CBI(5),
    CBI7  => CBI(6),
    CBI8  => CBI(7),
    CBI9  => CBI(8),
    CBI10 => CBI(9),
    CBI11 => CBI(10),
    CBI12 => CBI(11),
    CBI13 => CBI(12),
    CBI14 => CBI(13),
    CBI15 => CBI(14),
    CBI16 => CBI(15),
    CBI17 => CBI(16),
    CBI18 => CBI(17),

    CBO1  => CBO(0),
    CBO2  => CBO(1),
    CBO3  => CBO(2),
    CBO4  => CBO(3),
    CBO5  => CBO(4),
    CBO6  => CBO(5),
    CBO7  => CBO(6),
    CBO8  => CBO(7),
    CBO9  => CBO(8),
    CBO10 => CBO(9),
    CBO11 => CBO(10),
    CBO12 => CBO(11),
    CBO13 => CBO(12),
    CBO14 => CBO(13),
    CBO15 => CBO(14),
    CBO16 => CBO(15),
    CBO17 => CBO(16),
    CBO18 => CBO(17),

    CCI   => CCI,
    CCO   => CCO,
    CI    => CI,
    CK    => CK,
    CO    => CO,
    CO37  => CO37,
    CO57  => CO57,

    CZI1  => CZI(0),
    CZI2  => CZI(1),
    CZI3  => CZI(2),
    CZI4  => CZI(3),
    CZI5  => CZI(4),
    CZI6  => CZI(5),
    CZI7  => CZI(6),
    CZI8  => CZI(7),
    CZI9  => CZI(8),
    CZI10 => CZI(9),
    CZI11 => CZI(10),
    CZI12 => CZI(11),
    CZI13 => CZI(12),
    CZI14 => CZI(13),
    CZI15 => CZI(14),
    CZI16 => CZI(15),
    CZI17 => CZI(16),
    CZI18 => CZI(17),
    CZI19 => CZI(18),
    CZI20 => CZI(19),
    CZI21 => CZI(20),
    CZI22 => CZI(21),
    CZI23 => CZI(22),
    CZI24 => CZI(23),
    CZI25 => CZI(24),
    CZI26 => CZI(25),
    CZI27 => CZI(26),
    CZI28 => CZI(27),
    CZI29 => CZI(28),
    CZI30 => CZI(29),
    CZI31 => CZI(30),
    CZI32 => CZI(31),
    CZI33 => CZI(32),
    CZI34 => CZI(33),
    CZI35 => CZI(34),
    CZI36 => CZI(35),
    CZI37 => CZI(36),
    CZI38 => CZI(37),
    CZI39 => CZI(38),
    CZI40 => CZI(39),
    CZI41 => CZI(40),
    CZI42 => CZI(41),
    CZI43 => CZI(42),
    CZI44 => CZI(43),
    CZI45 => CZI(44),
    CZI46 => CZI(45),
    CZI47 => CZI(46),
    CZI48 => CZI(47),
    CZI49 => CZI(48),
    CZI50 => CZI(49),
    CZI51 => CZI(50),
    CZI52 => CZI(51),
    CZI53 => CZI(52),
    CZI54 => CZI(53),
    CZI55 => CZI(54),
    CZI56 => CZI(55),

    CZO1  => CZO(0),
    CZO2  => CZO(1),
    CZO3  => CZO(2),
    CZO4  => CZO(3),
    CZO5  => CZO(4),
    CZO6  => CZO(5),
    CZO7  => CZO(6),
    CZO8  => CZO(7),
    CZO9  => CZO(8),
    CZO10 => CZO(9),
    CZO11 => CZO(10),
    CZO12 => CZO(11),
    CZO13 => CZO(12),
    CZO14 => CZO(13),
    CZO15 => CZO(14),
    CZO16 => CZO(15),
    CZO17 => CZO(16),
    CZO18 => CZO(17),
    CZO19 => CZO(18),
    CZO20 => CZO(19),
    CZO21 => CZO(20),
    CZO22 => CZO(21),
    CZO23 => CZO(22),
    CZO24 => CZO(23),
    CZO25 => CZO(24),
    CZO26 => CZO(25),
    CZO27 => CZO(26),
    CZO28 => CZO(27),
    CZO29 => CZO(28),
    CZO30 => CZO(29),
    CZO31 => CZO(30),
    CZO32 => CZO(31),
    CZO33 => CZO(32),
    CZO34 => CZO(33),
    CZO35 => CZO(34),
    CZO36 => CZO(35),
    CZO37 => CZO(36),
    CZO38 => CZO(37),
    CZO39 => CZO(38),
    CZO40 => CZO(39),
    CZO41 => CZO(40),
    CZO42 => CZO(41),
    CZO43 => CZO(42),
    CZO44 => CZO(43),
    CZO45 => CZO(44),
    CZO46 => CZO(45),
    CZO47 => CZO(46),
    CZO48 => CZO(47),
    CZO49 => CZO(48),
    CZO50 => CZO(49),
    CZO51 => CZO(50),
    CZO52 => CZO(51),
    CZO53 => CZO(52),
    CZO54 => CZO(53),
    CZO55 => CZO(54),
    CZO56 => CZO(55),

    D1    => D(0),
    D2    => D(1),
    D3    => D(2),
    D4    => D(3),
    D5    => D(4),
    D6    => D(5),
    D7    => D(6),
    D8    => D(7),
    D9    => D(8),
    D10   => D(9),
    D11   => D(10),
    D12   => D(11),
    D13   => D(12),
    D14   => D(13),
    D15   => D(14),
    D16   => D(15),
    D17   => D(16),
    D18   => D(17),

    OVF   => OVF,
    R     => R,
    RZ    => RZ,
    WE    => WE,

    Z1    => Z(0),
    Z2    => Z(1),
    Z3    => Z(2),
    Z4    => Z(3),
    Z5    => Z(4),
    Z6    => Z(5),
    Z7    => Z(6),
    Z8    => Z(7),
    Z9    => Z(8),
    Z10   => Z(9),
    Z11   => Z(10),
    Z12   => Z(11),
    Z13   => Z(12),
    Z14   => Z(13),
    Z15   => Z(14),
    Z16   => Z(15),
    Z17   => Z(16),
    Z18   => Z(17),
    Z19   => Z(18),
    Z20   => Z(19),
    Z21   => Z(20),
    Z22   => Z(21),
    Z23   => Z(22),
    Z24   => Z(23),
    Z25   => Z(24),
    Z26   => Z(25),
    Z27   => Z(26),
    Z28   => Z(27),
    Z29   => Z(28),
    Z30   => Z(29),
    Z31   => Z(30),
    Z32   => Z(31),
    Z33   => Z(32),
    Z34   => Z(33),
    Z35   => Z(34),
    Z36   => Z(35),
    Z37   => Z(36),
    Z38   => Z(37),
    Z39   => Z(38),
    Z40   => Z(39),
    Z41   => Z(40),
    Z42   => Z(41),
    Z43   => Z(42),
    Z44   => Z(43),
    Z45   => Z(44),
    Z46   => Z(45),
    Z47   => Z(46),
    Z48   => Z(47),
    Z49   => Z(48),
    Z50   => Z(49),
    Z51   => Z(50),
    Z52   => Z(51),
    Z53   => Z(52),
    Z54   => Z(53),
    Z55   => Z(54),
    Z56   => Z(55)
);

end NX_ARCH;
-- #}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_L_SPLIT definition                                                          2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_signed.ALL;

entity NX_DSP_L_SPLIT is
generic (
-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
------------------------------------------------------------------------- 
   SIGNED_MODE          : bit                    := '0';
   PRE_ADDER_OP         : bit                    := '0';       -- '0' = Additon, '1' = Subraction
   MUX_A                : bit                    := '0';       -- '0' = A input, '1' = CAI input
   MUX_B                : bit                    := '0';       -- '0' = B input, '1' = CBI input
   MUX_P                : bit                    := '0';       -- '0' for PRE_ADDER, '0' for B input
   MUX_X                : bit_vector(1 downto 0) := B"00";     -- Select X operand   "00" = C,
                                                               --                    "01" = CZI,
                                                               --                    "11" = SHFT(CZI) & C(11:0),
                                                               --                    "10" Select Z feedback
   MUX_Y                : bit                    := '0';       -- '0' Select MULT output, '1' for (B & A)
   MUX_CI               : bit                    := '0';       -- Select fabric input (not cascade)
   MUX_Z                : bit                    := '0';       -- Select ALU output
                                                               -- (not ALU input operand coming from PR_Y)

   Z_FEEDBACK_SHL12     : bit                    := '0';       -- '0' for No shift, '1' for 12-bit left shift
   ENABLE_SATURATION    : bit                    := '0';       -- '0' for Disable,  '1' for Enable
   SATURATION_RANK      : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB
                                                               --        on Z and CZO result
                                                               --(to define saturation and overflow)

   ALU_DYNAMIC_OP       : bit                    := '0';       -- '0' for Static,
                                                               -- '1' for Dynamic
                                                               -- (D6 ... D1 is not used for dynamic operation)
   CO_SEL               : bit                    := '0';       -- '0' for C0 = ALU(36), '1' for CO = ALU(48)

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
-------------------------------------------------------------------------
   PR_A_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on A input
   PR_A_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output
   PR_B_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on B input
   PR_B_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output

   PR_C_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_D_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_CI_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_P_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
   PR_X_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_Y_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

   PR_MULT_MUX             : bit                    := '0';   -- No pipe reg  -- Register inside MULT
   PR_ALU_MUX              : bit                    := '0';   -- No pipe reg  -- Register inside ALU
   PR_Z_MUX                : bit                    := '0';   -- Registered output

   PR_CO_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_OV_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
-------------------------------------------------------------------------
   ENABLE_PR_A_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_B_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_C_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_D_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CI_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_P_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_X_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Y_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_MULT_RST      : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_ALU_RST       : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Z_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CO_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_OV_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 

-------------------------------------------------------------------------
-- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
-------------------------------------------------------------------------
   ALU_OP                  : bit_vector(5 downto 0) := B"000000"; -- Addition = "000000", Subtract = "001010"
   ALU_MUX                 : bit                    := '0'        -- '0' for Don't swap ALU operands,
                                                                  -- '1' for ALU Swap operands
    );
port(
   CK   : IN  std_logic;
   R    : IN  std_logic;
   RZ   : IN  std_logic;
   WE   : IN  std_logic;

   CI   : IN  std_logic;     -- cy_i
   A    : IN  std_logic_vector(23 downto 0);
   B    : IN  std_logic_vector(17 downto 0);
   C    : IN  std_logic_vector(35 downto 0);
   D    : IN  std_logic_vector(17 downto 0);
   CAI  : IN  std_logic_vector(23 downto 0);
   CBI  : IN  std_logic_vector(17 downto 0);
   CZI  : IN  std_logic_vector(55 downto 0);
   CCI  : IN  std_logic;  -- ccy_i

   Z    : out  std_logic_vector(55 downto 0);
   CO   : OUT  std_logic;  -- cy_o
   CO36 : OUT  std_logic;  -- cy36_o
   CO56 : OUT  std_logic;  -- cy56_o
   OVF  : OUT  std_logic;
   CAO  : OUT  std_logic_vector(23 downto 0);
   CBO  : OUT  std_logic_vector(17 downto 0);
   CZO  : OUT  std_logic_vector(55 downto 0);
   CCO  : OUT  std_logic  -- ccy_o
  );
end NX_DSP_L_SPLIT;

-- architecture NX_RTL of NX_DSP_L_SPLIT#{{{#
architecture NX_RTL of NX_DSP_L_SPLIT is

----------------------------------------------------------
-- Internal signals to be mapped to the NX_DSP_L component
----------------------------------------------------------
signal A1         : std_logic := '0';
signal A2         : std_logic := '0';
signal A3         : std_logic := '0';
signal A4         : std_logic := '0';
signal A5         : std_logic := '0';
signal A6         : std_logic := '0';
signal A7         : std_logic := '0';
signal A8         : std_logic := '0';
signal A9         : std_logic := '0';
signal A10        : std_logic := '0';
signal A11        : std_logic := '0';
signal A12        : std_logic := '0';
signal A13        : std_logic := '0';
signal A14        : std_logic := '0';
signal A15        : std_logic := '0';
signal A16        : std_logic := '0';
signal A17        : std_logic := '0';
signal A18        : std_logic := '0';
signal A19        : std_logic := '0';
signal A20        : std_logic := '0';
signal A21        : std_logic := '0';
signal A22        : std_logic := '0';
signal A23        : std_logic := '0';
signal A24        : std_logic := '0';

signal B1         : std_logic := '0';
signal B2         : std_logic := '0';
signal B3         : std_logic := '0';
signal B4         : std_logic := '0';
signal B5         : std_logic := '0';
signal B6         : std_logic := '0';
signal B7         : std_logic := '0';
signal B8         : std_logic := '0';
signal B9         : std_logic := '0';
signal B10        : std_logic := '0';
signal B11        : std_logic := '0';
signal B12        : std_logic := '0';
signal B13        : std_logic := '0';
signal B14        : std_logic := '0';
signal B15        : std_logic := '0';
signal B16        : std_logic := '0';
signal B17        : std_logic := '0';
signal B18        : std_logic := '0';
         
signal C1         : std_logic := '0';
signal C2         : std_logic := '0';
signal C3         : std_logic := '0';
signal C4         : std_logic := '0';
signal C5         : std_logic := '0';
signal C6         : std_logic := '0';
signal C7         : std_logic := '0';
signal C8         : std_logic := '0';
signal C9         : std_logic := '0';
signal C10        : std_logic := '0';
signal C11        : std_logic := '0';
signal C12        : std_logic := '0';
signal C13        : std_logic := '0';
signal C14        : std_logic := '0';
signal C15        : std_logic := '0';
signal C16        : std_logic := '0';
signal C17        : std_logic := '0';
signal C18        : std_logic := '0';
signal C19        : std_logic := '0';
signal C20        : std_logic := '0';
signal C21        : std_logic := '0';
signal C22        : std_logic := '0';
signal C23        : std_logic := '0';
signal C24        : std_logic := '0';
signal C25        : std_logic := '0';
signal C26        : std_logic := '0';
signal C27        : std_logic := '0';
signal C28        : std_logic := '0';
signal C29        : std_logic := '0';
signal C30        : std_logic := '0';
signal C31        : std_logic := '0';
signal C32        : std_logic := '0';
signal C33        : std_logic := '0';
signal C34        : std_logic := '0';
signal C35        : std_logic := '0';
signal C36        : std_logic := '0';

signal CAI1       : std_logic := '0';
signal CAI2       : std_logic := '0';
signal CAI3       : std_logic := '0';
signal CAI4       : std_logic := '0';
signal CAI5       : std_logic := '0';
signal CAI6       : std_logic := '0';
signal CAI7       : std_logic := '0';
signal CAI8       : std_logic := '0';
signal CAI9       : std_logic := '0';
signal CAI10      : std_logic := '0';
signal CAI11      : std_logic := '0';
signal CAI12      : std_logic := '0';
signal CAI13      : std_logic := '0';
signal CAI14      : std_logic := '0';
signal CAI15      : std_logic := '0';
signal CAI16      : std_logic := '0';
signal CAI17      : std_logic := '0';
signal CAI18      : std_logic := '0';
signal CAI19      : std_logic := '0';
signal CAI20      : std_logic := '0';
signal CAI21      : std_logic := '0';
signal CAI22      : std_logic := '0';
signal CAI23      : std_logic := '0';
signal CAI24      : std_logic := '0';

signal CAO1       : std_logic := '0';
signal CAO2       : std_logic := '0';
signal CAO3       : std_logic := '0';
signal CAO4       : std_logic := '0';
signal CAO5       : std_logic := '0';
signal CAO6       : std_logic := '0';
signal CAO7       : std_logic := '0';
signal CAO8       : std_logic := '0';
signal CAO9       : std_logic := '0';
signal CAO10      : std_logic := '0';
signal CAO11      : std_logic := '0';
signal CAO12      : std_logic := '0';
signal CAO13      : std_logic := '0';
signal CAO14      : std_logic := '0';
signal CAO15      : std_logic := '0';
signal CAO16      : std_logic := '0';
signal CAO17      : std_logic := '0';
signal CAO18      : std_logic := '0';
signal CAO19      : std_logic := '0';
signal CAO20      : std_logic := '0';
signal CAO21      : std_logic := '0';
signal CAO22      : std_logic := '0';
signal CAO23      : std_logic := '0';
signal CAO24      : std_logic := '0';

signal CBI1       : std_logic := '0';
signal CBI2       : std_logic := '0';
signal CBI3       : std_logic := '0';
signal CBI4       : std_logic := '0';
signal CBI5       : std_logic := '0';
signal CBI6       : std_logic := '0';
signal CBI7       : std_logic := '0';
signal CBI8       : std_logic := '0';
signal CBI9       : std_logic := '0';
signal CBI10      : std_logic := '0';
signal CBI11      : std_logic := '0';
signal CBI12      : std_logic := '0';
signal CBI13      : std_logic := '0';
signal CBI14      : std_logic := '0';
signal CBI15      : std_logic := '0';
signal CBI16      : std_logic := '0';
signal CBI17      : std_logic := '0';
signal CBI18      : std_logic := '0';

signal CBO1       : std_logic := '0';
signal CBO2       : std_logic := '0';
signal CBO3       : std_logic := '0';
signal CBO4       : std_logic := '0';
signal CBO5       : std_logic := '0';
signal CBO6       : std_logic := '0';
signal CBO7       : std_logic := '0';
signal CBO8       : std_logic := '0';
signal CBO9       : std_logic := '0';
signal CBO10      : std_logic := '0';
signal CBO11      : std_logic := '0';
signal CBO12      : std_logic := '0';
signal CBO13      : std_logic := '0';
signal CBO14      : std_logic := '0';
signal CBO15      : std_logic := '0';
signal CBO16      : std_logic := '0';
signal CBO17      : std_logic := '0';
signal CBO18      : std_logic := '0';

signal CO37       : std_logic := '0';
signal CO57       : std_logic := '0';

signal CZI1       : std_logic := '0';
signal CZI2       : std_logic := '0';
signal CZI3       : std_logic := '0';
signal CZI4       : std_logic := '0';
signal CZI5       : std_logic := '0';
signal CZI6       : std_logic := '0';
signal CZI7       : std_logic := '0';
signal CZI8       : std_logic := '0';
signal CZI9       : std_logic := '0';
signal CZI10      : std_logic := '0';
signal CZI11      : std_logic := '0';
signal CZI12      : std_logic := '0';
signal CZI13      : std_logic := '0';
signal CZI14      : std_logic := '0';
signal CZI15      : std_logic := '0';
signal CZI16      : std_logic := '0';
signal CZI17      : std_logic := '0';
signal CZI18      : std_logic := '0';
signal CZI19      : std_logic := '0';
signal CZI20      : std_logic := '0';
signal CZI21      : std_logic := '0';
signal CZI22      : std_logic := '0';
signal CZI23      : std_logic := '0';
signal CZI24      : std_logic := '0';
signal CZI25      : std_logic := '0';
signal CZI26      : std_logic := '0';
signal CZI27      : std_logic := '0';
signal CZI28      : std_logic := '0';
signal CZI29      : std_logic := '0';
signal CZI30      : std_logic := '0';
signal CZI31      : std_logic := '0';
signal CZI32      : std_logic := '0';
signal CZI33      : std_logic := '0';
signal CZI34      : std_logic := '0';
signal CZI35      : std_logic := '0';
signal CZI36      : std_logic := '0';
signal CZI37      : std_logic := '0';
signal CZI38      : std_logic := '0';
signal CZI39      : std_logic := '0';
signal CZI40      : std_logic := '0';
signal CZI41      : std_logic := '0';
signal CZI42      : std_logic := '0';
signal CZI43      : std_logic := '0';
signal CZI44      : std_logic := '0';
signal CZI45      : std_logic := '0';
signal CZI46      : std_logic := '0';
signal CZI47      : std_logic := '0';
signal CZI48      : std_logic := '0';
signal CZI49      : std_logic := '0';
signal CZI50      : std_logic := '0';
signal CZI51      : std_logic := '0';
signal CZI52      : std_logic := '0';
signal CZI53      : std_logic := '0';
signal CZI54      : std_logic := '0';
signal CZI55      : std_logic := '0';
signal CZI56      : std_logic := '0';

signal CZO1       : std_logic := '0';
signal CZO2       : std_logic := '0';
signal CZO3       : std_logic := '0';
signal CZO4       : std_logic := '0';
signal CZO5       : std_logic := '0';
signal CZO6       : std_logic := '0';
signal CZO7       : std_logic := '0';
signal CZO8       : std_logic := '0';
signal CZO9       : std_logic := '0';
signal CZO10      : std_logic := '0';
signal CZO11      : std_logic := '0';
signal CZO12      : std_logic := '0';
signal CZO13      : std_logic := '0';
signal CZO14      : std_logic := '0';
signal CZO15      : std_logic := '0';
signal CZO16      : std_logic := '0';
signal CZO17      : std_logic := '0';
signal CZO18      : std_logic := '0';
signal CZO19      : std_logic := '0';
signal CZO20      : std_logic := '0';
signal CZO21      : std_logic := '0';
signal CZO22      : std_logic := '0';
signal CZO23      : std_logic := '0';
signal CZO24      : std_logic := '0';
signal CZO25      : std_logic := '0';
signal CZO26      : std_logic := '0';
signal CZO27      : std_logic := '0';
signal CZO28      : std_logic := '0';
signal CZO29      : std_logic := '0';
signal CZO30      : std_logic := '0';
signal CZO31      : std_logic := '0';
signal CZO32      : std_logic := '0';
signal CZO33      : std_logic := '0';
signal CZO34      : std_logic := '0';
signal CZO35      : std_logic := '0';
signal CZO36      : std_logic := '0';
signal CZO37      : std_logic := '0';
signal CZO38      : std_logic := '0';
signal CZO39      : std_logic := '0';
signal CZO40      : std_logic := '0';
signal CZO41      : std_logic := '0';
signal CZO42      : std_logic := '0';
signal CZO43      : std_logic := '0';
signal CZO44      : std_logic := '0';
signal CZO45      : std_logic := '0';
signal CZO46      : std_logic := '0';
signal CZO47      : std_logic := '0';
signal CZO48      : std_logic := '0';
signal CZO49      : std_logic := '0';
signal CZO50      : std_logic := '0';
signal CZO51      : std_logic := '0';
signal CZO52      : std_logic := '0';
signal CZO53      : std_logic := '0';
signal CZO54      : std_logic := '0';
signal CZO55      : std_logic := '0';
signal CZO56      : std_logic := '0';

signal D1         : std_logic := '0';
signal D2         : std_logic := '0';
signal D3         : std_logic := '0';
signal D4         : std_logic := '0';
signal D5         : std_logic := '0';
signal D6         : std_logic := '0';
signal D7         : std_logic := '0';
signal D8         : std_logic := '0';
signal D9         : std_logic := '0';
signal D10        : std_logic := '0';
signal D11        : std_logic := '0';
signal D12        : std_logic := '0';
signal D13        : std_logic := '0';
signal D14        : std_logic := '0';
signal D15        : std_logic := '0';
signal D16        : std_logic := '0';
signal D17        : std_logic := '0';
signal D18        : std_logic := '0';

signal Z1         : std_logic := '0';
signal Z2         : std_logic := '0';
signal Z3         : std_logic := '0';
signal Z4         : std_logic := '0';
signal Z5         : std_logic := '0';
signal Z6         : std_logic := '0';
signal Z7         : std_logic := '0';
signal Z8         : std_logic := '0';
signal Z9         : std_logic := '0';
signal Z10        : std_logic := '0';
signal Z11        : std_logic := '0';
signal Z12        : std_logic := '0';
signal Z13        : std_logic := '0';
signal Z14        : std_logic := '0';
signal Z15        : std_logic := '0';
signal Z16        : std_logic := '0';
signal Z17        : std_logic := '0';
signal Z18        : std_logic := '0';
signal Z19        : std_logic := '0';
signal Z20        : std_logic := '0';
signal Z21        : std_logic := '0';
signal Z22        : std_logic := '0';
signal Z23        : std_logic := '0';
signal Z24        : std_logic := '0';
signal Z25        : std_logic := '0';
signal Z26        : std_logic := '0';
signal Z27        : std_logic := '0';
signal Z28        : std_logic := '0';
signal Z29        : std_logic := '0';
signal Z30        : std_logic := '0';
signal Z31        : std_logic := '0';
signal Z32        : std_logic := '0';
signal Z33        : std_logic := '0';
signal Z34        : std_logic := '0';
signal Z35        : std_logic := '0';
signal Z36        : std_logic := '0';
signal Z37        : std_logic := '0';
signal Z38        : std_logic := '0';
signal Z39        : std_logic := '0';
signal Z40        : std_logic := '0';
signal Z41        : std_logic := '0';
signal Z42        : std_logic := '0';
signal Z43        : std_logic := '0';
signal Z44        : std_logic := '0';
signal Z45        : std_logic := '0';
signal Z46        : std_logic := '0';
signal Z47        : std_logic := '0';
signal Z48        : std_logic := '0';
signal Z49        : std_logic := '0';
signal Z50        : std_logic := '0';
signal Z51        : std_logic := '0';
signal Z52        : std_logic := '0';
signal Z53        : std_logic := '0';
signal Z54        : std_logic := '0';
signal Z55        : std_logic := '0';


constant raw_config0_gen : bit_vector(19 downto 0)
    := CO_SEL & ALU_DYNAMIC_OP & SATURATION_RANK & ENABLE_SATURATION & Z_FEEDBACK_SHL12 & MUX_Z &
       MUX_CI & MUX_Y & MUX_X & MUX_P & MUX_B & MUX_A & PRE_ADDER_OP & SIGNED_MODE;

constant raw_config1_gen : bit_vector(18 downto 0)
    := PR_OV_MUX & PR_CO_MUX & PR_Z_MUX & PR_ALU_MUX & PR_MULT_MUX & PR_Y_MUX & PR_X_MUX &
       PR_P_MUX & PR_CI_MUX & PR_D_MUX & PR_C_MUX & PR_B_CASCADE_MUX & PR_B_MUX & PR_A_CASCADE_MUX &
       PR_A_MUX;

constant raw_config2_gen : bit_vector(12 downto 0)
    := ENABLE_PR_OV_RST & ENABLE_PR_CO_RST & ENABLE_PR_Z_RST & ENABLE_PR_ALU_RST &
       ENABLE_PR_MULT_RST & ENABLE_PR_Y_RST & ENABLE_PR_X_RST & ENABLE_PR_P_RST & ENABLE_PR_CI_RST &
       ENABLE_PR_D_RST & ENABLE_PR_C_RST & ENABLE_PR_B_RST & ENABLE_PR_A_RST;

constant raw_config3_gen : bit_vector(6 downto 0) := ALU_MUX & ALU_OP;


----------------------------------------------------------
-- NX_DSP_L declaration
----------------------------------------------------------
component NX_DSP_L
generic (
   std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
   raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
   raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
   raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
   raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
   );
port (
   A1         : in std_logic := '0';
   A2         : in std_logic := '0';
   A3         : in std_logic := '0';
   A4         : in std_logic := '0';
   A5         : in std_logic := '0';
   A6         : in std_logic := '0';
   A7         : in std_logic := '0';
   A8         : in std_logic := '0';
   A9         : in std_logic := '0';
   A10        : in std_logic := '0';
   A11        : in std_logic := '0';
   A12        : in std_logic := '0';
   A13        : in std_logic := '0';
   A14        : in std_logic := '0';
   A15        : in std_logic := '0';
   A16        : in std_logic := '0';
   A17        : in std_logic := '0';
   A18        : in std_logic := '0';
   A19        : in std_logic := '0';
   A20        : in std_logic := '0';
   A21        : in std_logic := '0';
   A22        : in std_logic := '0';
   A23        : in std_logic := '0';
   A24        : in std_logic := '0';

   B1         : in std_logic := '0';
   B2         : in std_logic := '0';
   B3         : in std_logic := '0';
   B4         : in std_logic := '0';
   B5         : in std_logic := '0';
   B6         : in std_logic := '0';
   B7         : in std_logic := '0';
   B8         : in std_logic := '0';
   B9         : in std_logic := '0';
   B10        : in std_logic := '0';
   B11        : in std_logic := '0';
   B12        : in std_logic := '0';
   B13        : in std_logic := '0';
   B14        : in std_logic := '0';
   B15        : in std_logic := '0';
   B16        : in std_logic := '0';
   B17        : in std_logic := '0';
   B18        : in std_logic := '0';

   C1         : in std_logic := '0';
   C2         : in std_logic := '0';
   C3         : in std_logic := '0';
   C4         : in std_logic := '0';
   C5         : in std_logic := '0';
   C6         : in std_logic := '0';
   C7         : in std_logic := '0';
   C8         : in std_logic := '0';
   C9         : in std_logic := '0';
   C10        : in std_logic := '0';
   C11        : in std_logic := '0';
   C12        : in std_logic := '0';
   C13        : in std_logic := '0';
   C14        : in std_logic := '0';
   C15        : in std_logic := '0';
   C16        : in std_logic := '0';
   C17        : in std_logic := '0';
   C18        : in std_logic := '0';
   C19        : in std_logic := '0';
   C20        : in std_logic := '0';
   C21        : in std_logic := '0';
   C22        : in std_logic := '0';
   C23        : in std_logic := '0';
   C24        : in std_logic := '0';
   C25        : in std_logic := '0';
   C26        : in std_logic := '0';
   C27        : in std_logic := '0';
   C28        : in std_logic := '0';
   C29        : in std_logic := '0';
   C30        : in std_logic := '0';
   C31        : in std_logic := '0';
   C32        : in std_logic := '0';
   C33        : in std_logic := '0';
   C34        : in std_logic := '0';
   C35        : in std_logic := '0';
   C36        : in std_logic := '0';

   CAI1       : in std_logic := '0';
   CAI2       : in std_logic := '0';
   CAI3       : in std_logic := '0';
   CAI4       : in std_logic := '0';
   CAI5       : in std_logic := '0';
   CAI6       : in std_logic := '0';
   CAI7       : in std_logic := '0';
   CAI8       : in std_logic := '0';
   CAI9       : in std_logic := '0';
   CAI10      : in std_logic := '0';
   CAI11      : in std_logic := '0';
   CAI12      : in std_logic := '0';
   CAI13      : in std_logic := '0';
   CAI14      : in std_logic := '0';
   CAI15      : in std_logic := '0';
   CAI16      : in std_logic := '0';
   CAI17      : in std_logic := '0';
   CAI18      : in std_logic := '0';
   CAI19      : in std_logic := '0';
   CAI20      : in std_logic := '0';
   CAI21      : in std_logic := '0';
   CAI22      : in std_logic := '0';
   CAI23      : in std_logic := '0';
   CAI24      : in std_logic := '0';

   CAO1       : out std_logic := '0';
   CAO2       : out std_logic := '0';
   CAO3       : out std_logic := '0';
   CAO4       : out std_logic := '0';
   CAO5       : out std_logic := '0';
   CAO6       : out std_logic := '0';
   CAO7       : out std_logic := '0';
   CAO8       : out std_logic := '0';
   CAO9       : out std_logic := '0';
   CAO10      : out std_logic := '0';
   CAO11      : out std_logic := '0';
   CAO12      : out std_logic := '0';
   CAO13      : out std_logic := '0';
   CAO14      : out std_logic := '0';
   CAO15      : out std_logic := '0';
   CAO16      : out std_logic := '0';
   CAO17      : out std_logic := '0';
   CAO18      : out std_logic := '0';
   CAO19      : out std_logic := '0';
   CAO20      : out std_logic := '0';
   CAO21      : out std_logic := '0';
   CAO22      : out std_logic := '0';
   CAO23      : out std_logic := '0';
   CAO24      : out std_logic := '0';

   CBI1       : in std_logic := '0';
   CBI2       : in std_logic := '0';
   CBI3       : in std_logic := '0';
   CBI4       : in std_logic := '0';
   CBI5       : in std_logic := '0';
   CBI6       : in std_logic := '0';
   CBI7       : in std_logic := '0';
   CBI8       : in std_logic := '0';
   CBI9       : in std_logic := '0';
   CBI10      : in std_logic := '0';
   CBI11      : in std_logic := '0';
   CBI12      : in std_logic := '0';
   CBI13      : in std_logic := '0';
   CBI14      : in std_logic := '0';
   CBI15      : in std_logic := '0';
   CBI16      : in std_logic := '0';
   CBI17      : in std_logic := '0';
   CBI18      : in std_logic := '0';

   CBO1       : out std_logic := '0';
   CBO2       : out std_logic := '0';
   CBO3       : out std_logic := '0';
   CBO4       : out std_logic := '0';
   CBO5       : out std_logic := '0';
   CBO6       : out std_logic := '0';
   CBO7       : out std_logic := '0';
   CBO8       : out std_logic := '0';
   CBO9       : out std_logic := '0';
   CBO10      : out std_logic := '0';
   CBO11      : out std_logic := '0';
   CBO12      : out std_logic := '0';
   CBO13      : out std_logic := '0';
   CBO14      : out std_logic := '0';
   CBO15      : out std_logic := '0';
   CBO16      : out std_logic := '0';
   CBO17      : out std_logic := '0';
   CBO18      : out std_logic := '0';

   CCI        : in std_logic := '0';
   CCO        : out std_logic := '0';
   CI         : in std_logic := '0';
   CK         : in std_logic := '0';
   CO         : out std_logic := '0';
   CO37       : out std_logic := '0';
   CO57       : out std_logic := '0';

   CZI1       : in std_logic := '0';
   CZI2       : in std_logic := '0';
   CZI3       : in std_logic := '0';
   CZI4       : in std_logic := '0';
   CZI5       : in std_logic := '0';
   CZI6       : in std_logic := '0';
   CZI7       : in std_logic := '0';
   CZI8       : in std_logic := '0';
   CZI9       : in std_logic := '0';
   CZI10      : in std_logic := '0';
   CZI11      : in std_logic := '0';
   CZI12      : in std_logic := '0';
   CZI13      : in std_logic := '0';
   CZI14      : in std_logic := '0';
   CZI15      : in std_logic := '0';
   CZI16      : in std_logic := '0';
   CZI17      : in std_logic := '0';
   CZI18      : in std_logic := '0';
   CZI19      : in std_logic := '0';
   CZI20      : in std_logic := '0';
   CZI21      : in std_logic := '0';
   CZI22      : in std_logic := '0';
   CZI23      : in std_logic := '0';
   CZI24      : in std_logic := '0';
   CZI25      : in std_logic := '0';
   CZI26      : in std_logic := '0';
   CZI27      : in std_logic := '0';
   CZI28      : in std_logic := '0';
   CZI29      : in std_logic := '0';
   CZI30      : in std_logic := '0';
   CZI31      : in std_logic := '0';
   CZI32      : in std_logic := '0';
   CZI33      : in std_logic := '0';
   CZI34      : in std_logic := '0';
   CZI35      : in std_logic := '0';
   CZI36      : in std_logic := '0';
   CZI37      : in std_logic := '0';
   CZI38      : in std_logic := '0';
   CZI39      : in std_logic := '0';
   CZI40      : in std_logic := '0';
   CZI41      : in std_logic := '0';
   CZI42      : in std_logic := '0';
   CZI43      : in std_logic := '0';
   CZI44      : in std_logic := '0';
   CZI45      : in std_logic := '0';
   CZI46      : in std_logic := '0';
   CZI47      : in std_logic := '0';
   CZI48      : in std_logic := '0';
   CZI49      : in std_logic := '0';
   CZI50      : in std_logic := '0';
   CZI51      : in std_logic := '0';
   CZI52      : in std_logic := '0';
   CZI53      : in std_logic := '0';
   CZI54      : in std_logic := '0';
   CZI55      : in std_logic := '0';
   CZI56      : in std_logic := '0';

   CZO1       : out std_logic := '0';
   CZO2       : out std_logic := '0';
   CZO3       : out std_logic := '0';
   CZO4       : out std_logic := '0';
   CZO5       : out std_logic := '0';
   CZO6       : out std_logic := '0';
   CZO7       : out std_logic := '0';
   CZO8       : out std_logic := '0';
   CZO9       : out std_logic := '0';
   CZO10      : out std_logic := '0';
   CZO11      : out std_logic := '0';
   CZO12      : out std_logic := '0';
   CZO13      : out std_logic := '0';
   CZO14      : out std_logic := '0';
   CZO15      : out std_logic := '0';
   CZO16      : out std_logic := '0';
   CZO17      : out std_logic := '0';
   CZO18      : out std_logic := '0';
   CZO19      : out std_logic := '0';
   CZO20      : out std_logic := '0';
   CZO21      : out std_logic := '0';
   CZO22      : out std_logic := '0';
   CZO23      : out std_logic := '0';
   CZO24      : out std_logic := '0';
   CZO25      : out std_logic := '0';
   CZO26      : out std_logic := '0';
   CZO27      : out std_logic := '0';
   CZO28      : out std_logic := '0';
   CZO29      : out std_logic := '0';
   CZO30      : out std_logic := '0';
   CZO31      : out std_logic := '0';
   CZO32      : out std_logic := '0';
   CZO33      : out std_logic := '0';
   CZO34      : out std_logic := '0';
   CZO35      : out std_logic := '0';
   CZO36      : out std_logic := '0';
   CZO37      : out std_logic := '0';
   CZO38      : out std_logic := '0';
   CZO39      : out std_logic := '0';
   CZO40      : out std_logic := '0';
   CZO41      : out std_logic := '0';
   CZO42      : out std_logic := '0';
   CZO43      : out std_logic := '0';
   CZO44      : out std_logic := '0';
   CZO45      : out std_logic := '0';
   CZO46      : out std_logic := '0';
   CZO47      : out std_logic := '0';
   CZO48      : out std_logic := '0';
   CZO49      : out std_logic := '0';
   CZO50      : out std_logic := '0';
   CZO51      : out std_logic := '0';
   CZO52      : out std_logic := '0';
   CZO53      : out std_logic := '0';
   CZO54      : out std_logic := '0';
   CZO55      : out std_logic := '0';
   CZO56      : out std_logic := '0';

   D1         : in std_logic := '0';
   D2         : in std_logic := '0';
   D3         : in std_logic := '0';
   D4         : in std_logic := '0';
   D5         : in std_logic := '0';
   D6         : in std_logic := '0';
   D7         : in std_logic := '0';
   D8         : in std_logic := '0';
   D9         : in std_logic := '0';
   D10        : in std_logic := '0';
   D11        : in std_logic := '0';
   D12        : in std_logic := '0';
   D13        : in std_logic := '0';
   D14        : in std_logic := '0';
   D15        : in std_logic := '0';
   D16        : in std_logic := '0';
   D17        : in std_logic := '0';
   D18        : in std_logic := '0';

   OVF        : out std_logic := '0';
   R          : in std_logic := '0';
   RZ         : in std_logic := '0';
   WE         : in std_logic := '0';

   Z1         : out std_logic := '0';
   Z2         : out std_logic := '0';
   Z3         : out std_logic := '0';
   Z4         : out std_logic := '0';
   Z5         : out std_logic := '0';
   Z6         : out std_logic := '0';
   Z7         : out std_logic := '0';
   Z8         : out std_logic := '0';
   Z9         : out std_logic := '0';
   Z10        : out std_logic := '0';
   Z11        : out std_logic := '0';
   Z12        : out std_logic := '0';
   Z13        : out std_logic := '0';
   Z14        : out std_logic := '0';
   Z15        : out std_logic := '0';
   Z16        : out std_logic := '0';
   Z17        : out std_logic := '0';
   Z18        : out std_logic := '0';
   Z19        : out std_logic := '0';
   Z20        : out std_logic := '0';
   Z21        : out std_logic := '0';
   Z22        : out std_logic := '0';
   Z23        : out std_logic := '0';
   Z24        : out std_logic := '0';
   Z25        : out std_logic := '0';
   Z26        : out std_logic := '0';
   Z27        : out std_logic := '0';
   Z28        : out std_logic := '0';
   Z29        : out std_logic := '0';
   Z30        : out std_logic := '0';
   Z31        : out std_logic := '0';
   Z32        : out std_logic := '0';
   Z33        : out std_logic := '0';
   Z34        : out std_logic := '0';
   Z35        : out std_logic := '0';
   Z36        : out std_logic := '0';
   Z37        : out std_logic := '0';
   Z38        : out std_logic := '0';
   Z39        : out std_logic := '0';
   Z40        : out std_logic := '0';
   Z41        : out std_logic := '0';
   Z42        : out std_logic := '0';
   Z43        : out std_logic := '0';
   Z44        : out std_logic := '0';
   Z45        : out std_logic := '0';
   Z46        : out std_logic := '0';
   Z47        : out std_logic := '0';
   Z48        : out std_logic := '0';
   Z49        : out std_logic := '0';
   Z50        : out std_logic := '0';
   Z51        : out std_logic := '0';
   Z52        : out std_logic := '0';
   Z53        : out std_logic := '0';
   Z54        : out std_logic := '0';
   Z55        : out std_logic := '0';
   Z56        : out std_logic := '0'
   );
end component;

begin

----------------------------------------------------------
-- Instantiation the NX_DSP_L component
----------------------------------------------------------
DSP_INST : NX_DSP_L
generic map (
   std_mode    => "", -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
   raw_config0 => raw_config0_gen, -- MODE and MUXes
   raw_config1 => raw_config1_gen, -- Pipeline Registers
   raw_config2 => raw_config2_gen, -- Reset Enable for internal registers
   raw_config3 => raw_config3_gen   -- ALU modes
   )
port map (
   A1         => A(0),
   A2         => A(1),
   A3         => A(2),
   A4         => A(3),
   A5         => A(4),
   A6         => A(5),
   A7         => A(6),
   A8         => A(7),
   A9         => A(8),
   A10        => A(9),
   A11        => A(10),
   A12        => A(11),
   A13        => A(12),
   A14        => A(13),
   A15        => A(14),
   A16        => A(15),
   A17        => A(16),
   A18        => A(17),
   A19        => A(18),
   A20        => A(19),
   A21        => A(20),
   A22        => A(21),
   A23        => A(22),
   A24        => A(23),
         
   B1         => B(0),
   B2         => B(1),
   B3         => B(2),
   B4         => B(3),
   B5         => B(4),
   B6         => B(5),
   B7         => B(6),
   B8         => B(7),
   B9         => B(8),
   B10        => B(9),
   B11        => B(10),
   B12        => B(11),
   B13        => B(12),
   B14        => B(13),
   B15        => B(14),
   B16        => B(15),
   B17        => B(16),
   B18        => B(17),
        
   C1         => C(0),
   C2         => C(1),
   C3         => C(2),
   C4         => C(3),
   C5         => C(4),
   C6         => C(5),
   C7         => C(6),
   C8         => C(7),
   C9         => C(8),
   C10        => C(9),
   C11        => C(10),
   C12        => C(11),
   C13        => C(12),
   C14        => C(13),
   C15        => C(14),
   C16        => C(15),
   C17        => C(16),
   C18        => C(17),
   C19        => C(18),
   C20        => C(19),
   C21        => C(20),
   C22        => C(21),
   C23        => C(22),
   C24        => C(23),
   C25        => C(24),
   C26        => C(25),
   C27        => C(26),
   C28        => C(27),
   C29        => C(28),
   C30        => C(29),
   C31        => C(30),
   C32        => C(31),
   C33        => C(32),
   C34        => C(33),
   C35        => C(34),
   C36        => C(35),

   CAI1       => CAI(0),
   CAI2       => CAI(1),
   CAI3       => CAI(2),
   CAI4       => CAI(3),
   CAI5       => CAI(4),
   CAI6       => CAI(5),
   CAI7       => CAI(6),
   CAI8       => CAI(7),
   CAI9       => CAI(8),
   CAI10      => CAI(9),
   CAI11      => CAI(10),
   CAI12      => CAI(11),
   CAI13      => CAI(12),
   CAI14      => CAI(13),
   CAI15      => CAI(14),
   CAI16      => CAI(15),
   CAI17      => CAI(16),
   CAI18      => CAI(17),
   CAI19      => CAI(18),
   CAI20      => CAI(19),
   CAI21      => CAI(20),
   CAI22      => CAI(21),
   CAI23      => CAI(22),
   CAI24      => CAI(23),

   CAO1       => CAO(0),
   CAO2       => CAO(1),
   CAO3       => CAO(2),
   CAO4       => CAO(3),
   CAO5       => CAO(4),
   CAO6       => CAO(5),
   CAO7       => CAO(6),
   CAO8       => CAO(7),
   CAO9       => CAO(8),
   CAO10      => CAO(9),
   CAO11      => CAO(10),
   CAO12      => CAO(11),
   CAO13      => CAO(12),
   CAO14      => CAO(13),
   CAO15      => CAO(14),
   CAO16      => CAO(15),
   CAO17      => CAO(16),
   CAO18      => CAO(17),
   CAO19      => CAO(18),
   CAO20      => CAO(19),
   CAO21      => CAO(20),
   CAO22      => CAO(21),
   CAO23      => CAO(22),
   CAO24      => CAO(23),

   CBI1       => CBI(0),
   CBI2       => CBI(1),
   CBI3       => CBI(2),
   CBI4       => CBI(3),
   CBI5       => CBI(4),
   CBI6       => CBI(5),
   CBI7       => CBI(6),
   CBI8       => CBI(7),
   CBI9       => CBI(8),
   CBI10      => CBI(9),
   CBI11      => CBI(10),
   CBI12      => CBI(11),
   CBI13      => CBI(12),
   CBI14      => CBI(13),
   CBI15      => CBI(14),
   CBI16      => CBI(15),
   CBI17      => CBI(16),
   CBI18      => CBI(17),

   CBO1       => CBO(0),
   CBO2       => CBO(1),
   CBO3       => CBO(2),
   CBO4       => CBO(3),
   CBO5       => CBO(4),
   CBO6       => CBO(5),
   CBO7       => CBO(6),
   CBO8       => CBO(7),
   CBO9       => CBO(8),
   CBO10      => CBO(9),
   CBO11      => CBO(10),
   CBO12      => CBO(11),
   CBO13      => CBO(12),
   CBO14      => CBO(13),
   CBO15      => CBO(14),
   CBO16      => CBO(15),
   CBO17      => CBO(16),
   CBO18      => CBO(17),

   CCI        => CCI,
   CCO        => CCO,
   CI         => CI,
   CK         => CK,
   CO         => CO,
   CO37       => CO36,
   CO57       => CO56,

   CZI1       => CZI(0),
   CZI2       => CZI(1),
   CZI3       => CZI(2),
   CZI4       => CZI(3),
   CZI5       => CZI(4),
   CZI6       => CZI(5),
   CZI7       => CZI(6),
   CZI8       => CZI(7),
   CZI9       => CZI(8),
   CZI10      => CZI(9),
   CZI11      => CZI(10),
   CZI12      => CZI(11),
   CZI13      => CZI(12),
   CZI14      => CZI(13),
   CZI15      => CZI(14),
   CZI16      => CZI(15),
   CZI17      => CZI(16),
   CZI18      => CZI(17),
   CZI19      => CZI(18),
   CZI20      => CZI(19),
   CZI21      => CZI(20),
   CZI22      => CZI(21),
   CZI23      => CZI(22),
   CZI24      => CZI(23),
   CZI25      => CZI(24),
   CZI26      => CZI(25),
   CZI27      => CZI(26),
   CZI28      => CZI(27),
   CZI29      => CZI(28),
   CZI30      => CZI(29),
   CZI31      => CZI(30),
   CZI32      => CZI(31),
   CZI33      => CZI(32),
   CZI34      => CZI(33),
   CZI35      => CZI(34),
   CZI36      => CZI(35),
   CZI37      => CZI(36),
   CZI38      => CZI(37),
   CZI39      => CZI(38),
   CZI40      => CZI(39),
   CZI41      => CZI(40),
   CZI42      => CZI(41),
   CZI43      => CZI(42),
   CZI44      => CZI(43),
   CZI45      => CZI(44),
   CZI46      => CZI(45),
   CZI47      => CZI(46),
   CZI48      => CZI(47),
   CZI49      => CZI(48),
   CZI50      => CZI(49),
   CZI51      => CZI(50),
   CZI52      => CZI(51),
   CZI53      => CZI(52),
   CZI54      => CZI(53),
   CZI55      => CZI(54),
   CZI56      => CZI(55),

   CZO1       => CZO(0),
   CZO2       => CZO(1),
   CZO3       => CZO(2),
   CZO4       => CZO(3),
   CZO5       => CZO(4),
   CZO6       => CZO(5),
   CZO7       => CZO(6),
   CZO8       => CZO(7),
   CZO9       => CZO(8),
   CZO10      => CZO(9),
   CZO11      => CZO(10),
   CZO12      => CZO(11),
   CZO13      => CZO(12),
   CZO14      => CZO(13),
   CZO15      => CZO(14),
   CZO16      => CZO(15),
   CZO17      => CZO(16),
   CZO18      => CZO(17),
   CZO19      => CZO(18),
   CZO20      => CZO(19),
   CZO21      => CZO(20),
   CZO22      => CZO(21),
   CZO23      => CZO(22),
   CZO24      => CZO(23),
   CZO25      => CZO(24),
   CZO26      => CZO(25),
   CZO27      => CZO(26),
   CZO28      => CZO(27),
   CZO29      => CZO(28),
   CZO30      => CZO(29),
   CZO31      => CZO(30),
   CZO32      => CZO(31),
   CZO33      => CZO(32),
   CZO34      => CZO(33),
   CZO35      => CZO(34),
   CZO36      => CZO(35),
   CZO37      => CZO(36),
   CZO38      => CZO(37),
   CZO39      => CZO(38),
   CZO40      => CZO(39),
   CZO41      => CZO(40),
   CZO42      => CZO(41),
   CZO43      => CZO(42),
   CZO44      => CZO(43),
   CZO45      => CZO(44),
   CZO46      => CZO(45),
   CZO47      => CZO(46),
   CZO48      => CZO(47),
   CZO49      => CZO(48),
   CZO50      => CZO(49),
   CZO51      => CZO(50),
   CZO52      => CZO(51),
   CZO53      => CZO(52),
   CZO54      => CZO(53),
   CZO55      => CZO(54),
   CZO56      => CZO(55),

   D1         => D(0),
   D2         => D(1),
   D3         => D(2),
   D4         => D(3),
   D5         => D(4),
   D6         => D(5),
   D7         => D(6),
   D8         => D(7),
   D9         => D(8),
   D10        => D(9),
   D11        => D(10),
   D12        => D(11),
   D13        => D(12),
   D14        => D(13),
   D15        => D(14),
   D16        => D(15),
   D17        => D(16),
   D18        => D(17),

   OVF        => OVF,
   R          => R,
   RZ         => RZ,
   WE         => WE,

   Z1         => Z(0),
   Z2         => Z(1),
   Z3         => Z(2),
   Z4         => Z(3),
   Z5         => Z(4),
   Z6         => Z(5),
   Z7         => Z(6),
   Z8         => Z(7),
   Z9         => Z(8),
   Z10        => Z(9),
   Z11        => Z(10),
   Z12        => Z(11),
   Z13        => Z(12),
   Z14        => Z(13),
   Z15        => Z(14),
   Z16        => Z(15),
   Z17        => Z(16),
   Z18        => Z(17),
   Z19        => Z(18),
   Z20        => Z(19),
   Z21        => Z(20),
   Z22        => Z(21),
   Z23        => Z(22),
   Z24        => Z(23),
   Z25        => Z(24),
   Z26        => Z(25),
   Z27        => Z(26),
   Z28        => Z(27),
   Z29        => Z(28),
   Z30        => Z(29),
   Z31        => Z(30),
   Z32        => Z(31),
   Z33        => Z(32),
   Z34        => Z(33),
   Z35        => Z(34),
   Z36        => Z(35),
   Z37        => Z(36),
   Z38        => Z(37),
   Z39        => Z(38),
   Z40        => Z(39),
   Z41        => Z(40),
   Z42        => Z(41),
   Z43        => Z(42),
   Z44        => Z(43),
   Z45        => Z(44),
   Z46        => Z(45),
   Z47        => Z(46),
   Z48        => Z(47),
   Z49        => Z(48),
   Z50        => Z(49),
   Z51        => Z(50),
   Z52        => Z(51),
   Z53        => Z(52),
   Z54        => Z(53),
   Z55        => Z(54),
   Z56        => Z(55)
   );

end NX_RTL;
-- #}}}#
-- =================================================================================================
--   NX_DSP definition                                                                  2018/11/30
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DSP is
generic (
    std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO49  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end NX_DSP;

-- =================================================================================================
--   NX_DSP_WRAP definition                                                             2017/09/25
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity NX_DSP_WRAP is
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
);
port (
    A    : in  std_logic_vector(23 downto 0);
    B    : in  std_logic_vector(17 downto 0);
    C    : in  std_logic_vector(35 downto 0);

    CAI  : in  std_logic_vector(17 downto 0);
    CAO  : out std_logic_vector(17 downto 0);
    CBI  : in  std_logic_vector(17 downto 0);
    CBO  : out std_logic_vector(17 downto 0);

    CCI  : in  std_logic;
    CCO  : out std_logic;
    CI   : in  std_logic;
    CK   : in  std_logic;
    CO   : out std_logic;
    CO37 : out std_logic;
    CO49 : out std_logic;

    CZI  : in  std_logic_vector(55 downto 0);
    CZO  : out std_logic_vector(55 downto 0);

    D    : in  std_logic_vector(17 downto 0);

    OVF  : out std_logic;
    R    : in  std_logic;
    RZ   : in  std_logic;
    WE   : in  std_logic;

    Z    : out std_logic_vector(55 downto 0)
);
end NX_DSP_WRAP;

-- architecture NX_ARCH of NX_DSP_WRAP#{{{#
architecture NX_ARCH of NX_DSP_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_ARCH: architecture is "WRAPPER";

component NX_DSP
generic (
    std_mode    : string := "";
    raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";      -- MUX
    raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";       -- PRC
    raw_config2 : bit_vector(12 downto 0) := B"0000000000000";             -- PRR
    raw_config3 : bit_vector( 6 downto 0) := B"0000000"                    -- ALU
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    CO    : out std_logic;
    CO37  : out std_logic;
    CO49  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end component;

begin

dsp: NX_DSP generic map (
    std_mode    => std_mode,
    raw_config0 => raw_config0,
    raw_config1 => raw_config1,
    raw_config2 => raw_config2,
    raw_config3 => raw_config3)
port map (
    A1    => A(0),
    A2    => A(1),
    A3    => A(2),
    A4    => A(3),
    A5    => A(4),
    A6    => A(5),
    A7    => A(6),
    A8    => A(7),
    A9    => A(8),
    A10   => A(9),
    A11   => A(10),
    A12   => A(11),
    A13   => A(12),
    A14   => A(13),
    A15   => A(14),
    A16   => A(15),
    A17   => A(16),
    A18   => A(17),
    A19   => A(18),
    A20   => A(19),
    A21   => A(20),
    A22   => A(21),
    A23   => A(22),
    A24   => A(23),

    B1    => B(0),
    B2    => B(1),
    B3    => B(2),
    B4    => B(3),
    B5    => B(4),
    B6    => B(5),
    B7    => B(6),
    B8    => B(7),
    B9    => B(8),
    B10   => B(9),
    B11   => B(10),
    B12   => B(11),
    B13   => B(12),
    B14   => B(13),
    B15   => B(14),
    B16   => B(15),
    B17   => B(16),
    B18   => B(17),

    C1    => C(0),
    C2    => C(1),
    C3    => C(2),
    C4    => C(3),
    C5    => C(4),
    C6    => C(5),
    C7    => C(6),
    C8    => C(7),
    C9    => C(8),
    C10   => C(9),
    C11   => C(10),
    C12   => C(11),
    C13   => C(12),
    C14   => C(13),
    C15   => C(14),
    C16   => C(15),
    C17   => C(16),
    C18   => C(17),
    C19   => C(18),
    C20   => C(19),
    C21   => C(20),
    C22   => C(21),
    C23   => C(22),
    C24   => C(23),
    C25   => C(24),
    C26   => C(25),
    C27   => C(26),
    C28   => C(27),
    C29   => C(28),
    C30   => C(29),
    C31   => C(30),
    C32   => C(31),
    C33   => C(32),
    C34   => C(33),
    C35   => C(34),
    C36   => C(35),

    CAI1  => CAI(0),
    CAI2  => CAI(1),
    CAI3  => CAI(2),
    CAI4  => CAI(3),
    CAI5  => CAI(4),
    CAI6  => CAI(5),
    CAI7  => CAI(6),
    CAI8  => CAI(7),
    CAI9  => CAI(8),
    CAI10 => CAI(9),
    CAI11 => CAI(10),
    CAI12 => CAI(11),
    CAI13 => CAI(12),
    CAI14 => CAI(13),
    CAI15 => CAI(14),
    CAI16 => CAI(15),
    CAI17 => CAI(16),
    CAI18 => CAI(17),

    CAO1  => CAO(0),
    CAO2  => CAO(1),
    CAO3  => CAO(2),
    CAO4  => CAO(3),
    CAO5  => CAO(4),
    CAO6  => CAO(5),
    CAO7  => CAO(6),
    CAO8  => CAO(7),
    CAO9  => CAO(8),
    CAO10 => CAO(9),
    CAO11 => CAO(10),
    CAO12 => CAO(11),
    CAO13 => CAO(12),
    CAO14 => CAO(13),
    CAO15 => CAO(14),
    CAO16 => CAO(15),
    CAO17 => CAO(16),
    CAO18 => CAO(17),

    CBI1  => CBI(0),
    CBI2  => CBI(1),
    CBI3  => CBI(2),
    CBI4  => CBI(3),
    CBI5  => CBI(4),
    CBI6  => CBI(5),
    CBI7  => CBI(6),
    CBI8  => CBI(7),
    CBI9  => CBI(8),
    CBI10 => CBI(9),
    CBI11 => CBI(10),
    CBI12 => CBI(11),
    CBI13 => CBI(12),
    CBI14 => CBI(13),
    CBI15 => CBI(14),
    CBI16 => CBI(15),
    CBI17 => CBI(16),
    CBI18 => CBI(17),

    CBO1  => CBO(0),
    CBO2  => CBO(1),
    CBO3  => CBO(2),
    CBO4  => CBO(3),
    CBO5  => CBO(4),
    CBO6  => CBO(5),
    CBO7  => CBO(6),
    CBO8  => CBO(7),
    CBO9  => CBO(8),
    CBO10 => CBO(9),
    CBO11 => CBO(10),
    CBO12 => CBO(11),
    CBO13 => CBO(12),
    CBO14 => CBO(13),
    CBO15 => CBO(14),
    CBO16 => CBO(15),
    CBO17 => CBO(16),
    CBO18 => CBO(17),

    CCI   => CCI,
    CCO   => CCO,
    CI    => CI,
    CK    => CK,
    CO    => CO,
    CO37  => CO37,
    CO49  => CO49,

    CZI1  => CZI(0),
    CZI2  => CZI(1),
    CZI3  => CZI(2),
    CZI4  => CZI(3),
    CZI5  => CZI(4),
    CZI6  => CZI(5),
    CZI7  => CZI(6),
    CZI8  => CZI(7),
    CZI9  => CZI(8),
    CZI10 => CZI(9),
    CZI11 => CZI(10),
    CZI12 => CZI(11),
    CZI13 => CZI(12),
    CZI14 => CZI(13),
    CZI15 => CZI(14),
    CZI16 => CZI(15),
    CZI17 => CZI(16),
    CZI18 => CZI(17),
    CZI19 => CZI(18),
    CZI20 => CZI(19),
    CZI21 => CZI(20),
    CZI22 => CZI(21),
    CZI23 => CZI(22),
    CZI24 => CZI(23),
    CZI25 => CZI(24),
    CZI26 => CZI(25),
    CZI27 => CZI(26),
    CZI28 => CZI(27),
    CZI29 => CZI(28),
    CZI30 => CZI(29),
    CZI31 => CZI(30),
    CZI32 => CZI(31),
    CZI33 => CZI(32),
    CZI34 => CZI(33),
    CZI35 => CZI(34),
    CZI36 => CZI(35),
    CZI37 => CZI(36),
    CZI38 => CZI(37),
    CZI39 => CZI(38),
    CZI40 => CZI(39),
    CZI41 => CZI(40),
    CZI42 => CZI(41),
    CZI43 => CZI(42),
    CZI44 => CZI(43),
    CZI45 => CZI(44),
    CZI46 => CZI(45),
    CZI47 => CZI(46),
    CZI48 => CZI(47),
    CZI49 => CZI(48),
    CZI50 => CZI(49),
    CZI51 => CZI(50),
    CZI52 => CZI(51),
    CZI53 => CZI(52),
    CZI54 => CZI(53),
    CZI55 => CZI(54),
    CZI56 => CZI(55),

    CZO1  => CZO(0),
    CZO2  => CZO(1),
    CZO3  => CZO(2),
    CZO4  => CZO(3),
    CZO5  => CZO(4),
    CZO6  => CZO(5),
    CZO7  => CZO(6),
    CZO8  => CZO(7),
    CZO9  => CZO(8),
    CZO10 => CZO(9),
    CZO11 => CZO(10),
    CZO12 => CZO(11),
    CZO13 => CZO(12),
    CZO14 => CZO(13),
    CZO15 => CZO(14),
    CZO16 => CZO(15),
    CZO17 => CZO(16),
    CZO18 => CZO(17),
    CZO19 => CZO(18),
    CZO20 => CZO(19),
    CZO21 => CZO(20),
    CZO22 => CZO(21),
    CZO23 => CZO(22),
    CZO24 => CZO(23),
    CZO25 => CZO(24),
    CZO26 => CZO(25),
    CZO27 => CZO(26),
    CZO28 => CZO(27),
    CZO29 => CZO(28),
    CZO30 => CZO(29),
    CZO31 => CZO(30),
    CZO32 => CZO(31),
    CZO33 => CZO(32),
    CZO34 => CZO(33),
    CZO35 => CZO(34),
    CZO36 => CZO(35),
    CZO37 => CZO(36),
    CZO38 => CZO(37),
    CZO39 => CZO(38),
    CZO40 => CZO(39),
    CZO41 => CZO(40),
    CZO42 => CZO(41),
    CZO43 => CZO(42),
    CZO44 => CZO(43),
    CZO45 => CZO(44),
    CZO46 => CZO(45),
    CZO47 => CZO(46),
    CZO48 => CZO(47),
    CZO49 => CZO(48),
    CZO50 => CZO(49),
    CZO51 => CZO(50),
    CZO52 => CZO(51),
    CZO53 => CZO(52),
    CZO54 => CZO(53),
    CZO55 => CZO(54),
    CZO56 => CZO(55),

    D1    => D(0),
    D2    => D(1),
    D3    => D(2),
    D4    => D(3),
    D5    => D(4),
    D6    => D(5),
    D7    => D(6),
    D8    => D(7),
    D9    => D(8),
    D10   => D(9),
    D11   => D(10),
    D12   => D(11),
    D13   => D(12),
    D14   => D(13),
    D15   => D(14),
    D16   => D(15),
    D17   => D(16),
    D18   => D(17),

    OVF   => OVF,
    R     => R,
    RZ    => RZ,
    WE    => WE,

    Z1    => Z(0),
    Z2    => Z(1),
    Z3    => Z(2),
    Z4    => Z(3),
    Z5    => Z(4),
    Z6    => Z(5),
    Z7    => Z(6),
    Z8    => Z(7),
    Z9    => Z(8),
    Z10   => Z(9),
    Z11   => Z(10),
    Z12   => Z(11),
    Z13   => Z(12),
    Z14   => Z(13),
    Z15   => Z(14),
    Z16   => Z(15),
    Z17   => Z(16),
    Z18   => Z(17),
    Z19   => Z(18),
    Z20   => Z(19),
    Z21   => Z(20),
    Z22   => Z(21),
    Z23   => Z(22),
    Z24   => Z(23),
    Z25   => Z(24),
    Z26   => Z(25),
    Z27   => Z(26),
    Z28   => Z(27),
    Z29   => Z(28),
    Z30   => Z(29),
    Z31   => Z(30),
    Z32   => Z(31),
    Z33   => Z(32),
    Z34   => Z(33),
    Z35   => Z(34),
    Z36   => Z(35),
    Z37   => Z(36),
    Z38   => Z(37),
    Z39   => Z(38),
    Z40   => Z(39),
    Z41   => Z(40),
    Z42   => Z(41),
    Z43   => Z(42),
    Z44   => Z(43),
    Z45   => Z(44),
    Z46   => Z(45),
    Z47   => Z(46),
    Z48   => Z(47),
    Z49   => Z(48),
    Z50   => Z(49),
    Z51   => Z(50),
    Z52   => Z(51),
    Z53   => Z(52),
    Z54   => Z(53),
    Z55   => Z(54),
    Z56   => Z(55)
);

end NX_ARCH;
-- #}}}#

-- =================================================================================================
--   NX_DSP_SPLIT definition                                                             2017/09/25
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_signed.ALL;

entity NX_DSP_SPLIT is
generic (
-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
------------------------------------------------------------------------- 
   SIGNED_MODE          : bit                    := '0';
   PRE_ADDER_OP         : bit                    := '0';       -- '0' = Additon, '1' = Subraction
   MUX_A                : bit                    := '0';       -- '0' = A input, '1' = CAI input
   MUX_B                : bit                    := '0';       -- '0' = B input, '1' = CBI input
   MUX_P                : bit                    := '0';       -- '0' for PRE_ADDER, '0' for B input
   MUX_X                : bit_vector(1 downto 0) := B"00";     -- Select X operand   "00" = C,
                                                               --                    "01" = CZI,
                                                               --                    "11" = SHFT(CZI) & C(11:0),
                                                               --                    "10" Select Z feedback
   MUX_Y                : bit                    := '0';       -- '0' Select MULT output, '1' for (B & A)
   MUX_CI               : bit                    := '0';       -- Select fabric input (not cascade)
   MUX_Z                : bit                    := '0';       -- Select ALU output
                                                               -- (not ALU input operand coming from PR_Y)

   Z_FEEDBACK_SHL12     : bit                    := '0';       -- '0' for No shift, '1' for 12-bit left shift
   ENABLE_SATURATION    : bit                    := '0';       -- '0' for Disable,  '1' for Enable
   SATURATION_RANK      : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB
                                                               --        on Z and CZO result
                                                               --(to define saturation and overflow)

   ALU_DYNAMIC_OP       : bit                    := '0';       -- '0' for Static,
                                                               -- '1' for Dynamic
                                                               -- (D6 ... D1 is not used for dynamic operation)
   CO_SEL               : bit                    := '0';       -- '0' for C0 = ALU(36), '1' for CO = ALU(48)

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
-------------------------------------------------------------------------
   PR_A_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on A input
   PR_A_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output
   PR_B_MUX                : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        on B input
   PR_B_CASCADE_MUX        : bit_vector(1 downto 0) := B"00"; -- Number of pipe reg levels
                                                              --        for CAO output

   PR_C_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_D_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_CI_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_P_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
   PR_X_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_Y_MUX                : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

   PR_MULT_MUX             : bit                    := '0';   -- No pipe reg  -- Register inside MULT
   PR_ALU_MUX              : bit                    := '0';   -- No pipe reg  -- Register inside ALU
   PR_Z_MUX                : bit                    := '0';   -- Registered output

   PR_CO_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg
   PR_OV_MUX               : bit                    := '0';   -- '0' for No pipe reg, '1' for 1 pipe reg

-------------------------------------------------------------------------
-- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
-------------------------------------------------------------------------
   ENABLE_PR_A_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_B_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_C_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_D_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CI_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_P_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_X_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Y_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_MULT_RST      : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_ALU_RST       : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_Z_RST         : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_CO_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 
   ENABLE_PR_OV_RST        : bit                    := '0';   -- '0' for Disable, '1' for Enable 

-------------------------------------------------------------------------
-- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
-------------------------------------------------------------------------
   ALU_OP                  : bit_vector(5 downto 0) := B"000000"; -- Addition = "000000", Subtract = "001010"
   ALU_MUX                 : bit                    := '0'        -- '0' for Don't swap ALU operands,
                                                                  -- '1' for ALU Swap operands
    );
port(
   CK   : IN  std_logic;
   R    : IN  std_logic;
   RZ   : IN  std_logic;
   WE   : IN  std_logic;

   CI   : IN  std_logic;     -- cy_i
   A    : IN  std_logic_vector(23 downto 0);
   B    : IN  std_logic_vector(17 downto 0);
   C    : IN  std_logic_vector(35 downto 0);
   D    : IN  std_logic_vector(17 downto 0);
   CAI  : IN  std_logic_vector(17 downto 0);
   CBI  : IN  std_logic_vector(17 downto 0);
   CZI  : IN  std_logic_vector(55 downto 0);
   CCI  : IN  std_logic;  -- ccy_i

   Z    : out  std_logic_vector(55 downto 0);
   CO   : OUT  std_logic;  -- cy_o
   CO36 : OUT  std_logic;  -- cy36_o
   CO48 : OUT  std_logic;  -- cy48_o
   OVF  : OUT  std_logic;
   CAO  : OUT  std_logic_vector(17 downto 0);
   CBO  : OUT  std_logic_vector(17 downto 0);
   CZO  : OUT  std_logic_vector(55 downto 0);
   CCO  : OUT  std_logic  -- ccy_o
  );
end NX_DSP_SPLIT;

-- architecture NX_RTL of NX_DSP_SPLIT#{{{#
architecture NX_RTL of NX_DSP_SPLIT is

----------------------------------------------------------
-- Internal signals to be mapped to the NX_DSP component
----------------------------------------------------------
signal A1         : std_logic := '0';
signal A2         : std_logic := '0';
signal A3         : std_logic := '0';
signal A4         : std_logic := '0';
signal A5         : std_logic := '0';
signal A6         : std_logic := '0';
signal A7         : std_logic := '0';
signal A8         : std_logic := '0';
signal A9         : std_logic := '0';
signal A10        : std_logic := '0';
signal A11        : std_logic := '0';
signal A12        : std_logic := '0';
signal A13        : std_logic := '0';
signal A14        : std_logic := '0';
signal A15        : std_logic := '0';
signal A16        : std_logic := '0';
signal A17        : std_logic := '0';
signal A18        : std_logic := '0';
signal A19        : std_logic := '0';
signal A20        : std_logic := '0';
signal A21        : std_logic := '0';
signal A22        : std_logic := '0';
signal A23        : std_logic := '0';
signal A24        : std_logic := '0';

signal B1         : std_logic := '0';
signal B2         : std_logic := '0';
signal B3         : std_logic := '0';
signal B4         : std_logic := '0';
signal B5         : std_logic := '0';
signal B6         : std_logic := '0';
signal B7         : std_logic := '0';
signal B8         : std_logic := '0';
signal B9         : std_logic := '0';
signal B10        : std_logic := '0';
signal B11        : std_logic := '0';
signal B12        : std_logic := '0';
signal B13        : std_logic := '0';
signal B14        : std_logic := '0';
signal B15        : std_logic := '0';
signal B16        : std_logic := '0';
signal B17        : std_logic := '0';
signal B18        : std_logic := '0';
         
signal C1         : std_logic := '0';
signal C2         : std_logic := '0';
signal C3         : std_logic := '0';
signal C4         : std_logic := '0';
signal C5         : std_logic := '0';
signal C6         : std_logic := '0';
signal C7         : std_logic := '0';
signal C8         : std_logic := '0';
signal C9         : std_logic := '0';
signal C10        : std_logic := '0';
signal C11        : std_logic := '0';
signal C12        : std_logic := '0';
signal C13        : std_logic := '0';
signal C14        : std_logic := '0';
signal C15        : std_logic := '0';
signal C16        : std_logic := '0';
signal C17        : std_logic := '0';
signal C18        : std_logic := '0';
signal C19        : std_logic := '0';
signal C20        : std_logic := '0';
signal C21        : std_logic := '0';
signal C22        : std_logic := '0';
signal C23        : std_logic := '0';
signal C24        : std_logic := '0';
signal C25        : std_logic := '0';
signal C26        : std_logic := '0';
signal C27        : std_logic := '0';
signal C28        : std_logic := '0';
signal C29        : std_logic := '0';
signal C30        : std_logic := '0';
signal C31        : std_logic := '0';
signal C32        : std_logic := '0';
signal C33        : std_logic := '0';
signal C34        : std_logic := '0';
signal C35        : std_logic := '0';
signal C36        : std_logic := '0';

signal CAI1       : std_logic := '0';
signal CAI2       : std_logic := '0';
signal CAI3       : std_logic := '0';
signal CAI4       : std_logic := '0';
signal CAI5       : std_logic := '0';
signal CAI6       : std_logic := '0';
signal CAI7       : std_logic := '0';
signal CAI8       : std_logic := '0';
signal CAI9       : std_logic := '0';
signal CAI10      : std_logic := '0';
signal CAI11      : std_logic := '0';
signal CAI12      : std_logic := '0';
signal CAI13      : std_logic := '0';
signal CAI14      : std_logic := '0';
signal CAI15      : std_logic := '0';
signal CAI16      : std_logic := '0';
signal CAI17      : std_logic := '0';
signal CAI18      : std_logic := '0';

signal CAO1       : std_logic := '0';
signal CAO2       : std_logic := '0';
signal CAO3       : std_logic := '0';
signal CAO4       : std_logic := '0';
signal CAO5       : std_logic := '0';
signal CAO6       : std_logic := '0';
signal CAO7       : std_logic := '0';
signal CAO8       : std_logic := '0';
signal CAO9       : std_logic := '0';
signal CAO10      : std_logic := '0';
signal CAO11      : std_logic := '0';
signal CAO12      : std_logic := '0';
signal CAO13      : std_logic := '0';
signal CAO14      : std_logic := '0';
signal CAO15      : std_logic := '0';
signal CAO16      : std_logic := '0';
signal CAO17      : std_logic := '0';
signal CAO18      : std_logic := '0';

signal CBI1       : std_logic := '0';
signal CBI2       : std_logic := '0';
signal CBI3       : std_logic := '0';
signal CBI4       : std_logic := '0';
signal CBI5       : std_logic := '0';
signal CBI6       : std_logic := '0';
signal CBI7       : std_logic := '0';
signal CBI8       : std_logic := '0';
signal CBI9       : std_logic := '0';
signal CBI10      : std_logic := '0';
signal CBI11      : std_logic := '0';
signal CBI12      : std_logic := '0';
signal CBI13      : std_logic := '0';
signal CBI14      : std_logic := '0';
signal CBI15      : std_logic := '0';
signal CBI16      : std_logic := '0';
signal CBI17      : std_logic := '0';
signal CBI18      : std_logic := '0';

signal CBO1       : std_logic := '0';
signal CBO2       : std_logic := '0';
signal CBO3       : std_logic := '0';
signal CBO4       : std_logic := '0';
signal CBO5       : std_logic := '0';
signal CBO6       : std_logic := '0';
signal CBO7       : std_logic := '0';
signal CBO8       : std_logic := '0';
signal CBO9       : std_logic := '0';
signal CBO10      : std_logic := '0';
signal CBO11      : std_logic := '0';
signal CBO12      : std_logic := '0';
signal CBO13      : std_logic := '0';
signal CBO14      : std_logic := '0';
signal CBO15      : std_logic := '0';
signal CBO16      : std_logic := '0';
signal CBO17      : std_logic := '0';
signal CBO18      : std_logic := '0';

signal CO37       : std_logic := '0';
signal CO49       : std_logic := '0';

signal CZI1       : std_logic := '0';
signal CZI2       : std_logic := '0';
signal CZI3       : std_logic := '0';
signal CZI4       : std_logic := '0';
signal CZI5       : std_logic := '0';
signal CZI6       : std_logic := '0';
signal CZI7       : std_logic := '0';
signal CZI8       : std_logic := '0';
signal CZI9       : std_logic := '0';
signal CZI10      : std_logic := '0';
signal CZI11      : std_logic := '0';
signal CZI12      : std_logic := '0';
signal CZI13      : std_logic := '0';
signal CZI14      : std_logic := '0';
signal CZI15      : std_logic := '0';
signal CZI16      : std_logic := '0';
signal CZI17      : std_logic := '0';
signal CZI18      : std_logic := '0';
signal CZI19      : std_logic := '0';
signal CZI20      : std_logic := '0';
signal CZI21      : std_logic := '0';
signal CZI22      : std_logic := '0';
signal CZI23      : std_logic := '0';
signal CZI24      : std_logic := '0';
signal CZI25      : std_logic := '0';
signal CZI26      : std_logic := '0';
signal CZI27      : std_logic := '0';
signal CZI28      : std_logic := '0';
signal CZI29      : std_logic := '0';
signal CZI30      : std_logic := '0';
signal CZI31      : std_logic := '0';
signal CZI32      : std_logic := '0';
signal CZI33      : std_logic := '0';
signal CZI34      : std_logic := '0';
signal CZI35      : std_logic := '0';
signal CZI36      : std_logic := '0';
signal CZI37      : std_logic := '0';
signal CZI38      : std_logic := '0';
signal CZI39      : std_logic := '0';
signal CZI40      : std_logic := '0';
signal CZI41      : std_logic := '0';
signal CZI42      : std_logic := '0';
signal CZI43      : std_logic := '0';
signal CZI44      : std_logic := '0';
signal CZI45      : std_logic := '0';
signal CZI46      : std_logic := '0';
signal CZI47      : std_logic := '0';
signal CZI48      : std_logic := '0';
signal CZI49      : std_logic := '0';
signal CZI50      : std_logic := '0';
signal CZI51      : std_logic := '0';
signal CZI52      : std_logic := '0';
signal CZI53      : std_logic := '0';
signal CZI54      : std_logic := '0';
signal CZI55      : std_logic := '0';
signal CZI56      : std_logic := '0';

signal CZO1       : std_logic := '0';
signal CZO2       : std_logic := '0';
signal CZO3       : std_logic := '0';
signal CZO4       : std_logic := '0';
signal CZO5       : std_logic := '0';
signal CZO6       : std_logic := '0';
signal CZO7       : std_logic := '0';
signal CZO8       : std_logic := '0';
signal CZO9       : std_logic := '0';
signal CZO10      : std_logic := '0';
signal CZO11      : std_logic := '0';
signal CZO12      : std_logic := '0';
signal CZO13      : std_logic := '0';
signal CZO14      : std_logic := '0';
signal CZO15      : std_logic := '0';
signal CZO16      : std_logic := '0';
signal CZO17      : std_logic := '0';
signal CZO18      : std_logic := '0';
signal CZO19      : std_logic := '0';
signal CZO20      : std_logic := '0';
signal CZO21      : std_logic := '0';
signal CZO22      : std_logic := '0';
signal CZO23      : std_logic := '0';
signal CZO24      : std_logic := '0';
signal CZO25      : std_logic := '0';
signal CZO26      : std_logic := '0';
signal CZO27      : std_logic := '0';
signal CZO28      : std_logic := '0';
signal CZO29      : std_logic := '0';
signal CZO30      : std_logic := '0';
signal CZO31      : std_logic := '0';
signal CZO32      : std_logic := '0';
signal CZO33      : std_logic := '0';
signal CZO34      : std_logic := '0';
signal CZO35      : std_logic := '0';
signal CZO36      : std_logic := '0';
signal CZO37      : std_logic := '0';
signal CZO38      : std_logic := '0';
signal CZO39      : std_logic := '0';
signal CZO40      : std_logic := '0';
signal CZO41      : std_logic := '0';
signal CZO42      : std_logic := '0';
signal CZO43      : std_logic := '0';
signal CZO44      : std_logic := '0';
signal CZO45      : std_logic := '0';
signal CZO46      : std_logic := '0';
signal CZO47      : std_logic := '0';
signal CZO48      : std_logic := '0';
signal CZO49      : std_logic := '0';
signal CZO50      : std_logic := '0';
signal CZO51      : std_logic := '0';
signal CZO52      : std_logic := '0';
signal CZO53      : std_logic := '0';
signal CZO54      : std_logic := '0';
signal CZO55      : std_logic := '0';
signal CZO56      : std_logic := '0';

signal D1         : std_logic := '0';
signal D2         : std_logic := '0';
signal D3         : std_logic := '0';
signal D4         : std_logic := '0';
signal D5         : std_logic := '0';
signal D6         : std_logic := '0';
signal D7         : std_logic := '0';
signal D8         : std_logic := '0';
signal D9         : std_logic := '0';
signal D10        : std_logic := '0';
signal D11        : std_logic := '0';
signal D12        : std_logic := '0';
signal D13        : std_logic := '0';
signal D14        : std_logic := '0';
signal D15        : std_logic := '0';
signal D16        : std_logic := '0';
signal D17        : std_logic := '0';
signal D18        : std_logic := '0';

signal Z1         : std_logic := '0';
signal Z2         : std_logic := '0';
signal Z3         : std_logic := '0';
signal Z4         : std_logic := '0';
signal Z5         : std_logic := '0';
signal Z6         : std_logic := '0';
signal Z7         : std_logic := '0';
signal Z8         : std_logic := '0';
signal Z9         : std_logic := '0';
signal Z10        : std_logic := '0';
signal Z11        : std_logic := '0';
signal Z12        : std_logic := '0';
signal Z13        : std_logic := '0';
signal Z14        : std_logic := '0';
signal Z15        : std_logic := '0';
signal Z16        : std_logic := '0';
signal Z17        : std_logic := '0';
signal Z18        : std_logic := '0';
signal Z19        : std_logic := '0';
signal Z20        : std_logic := '0';
signal Z21        : std_logic := '0';
signal Z22        : std_logic := '0';
signal Z23        : std_logic := '0';
signal Z24        : std_logic := '0';
signal Z25        : std_logic := '0';
signal Z26        : std_logic := '0';
signal Z27        : std_logic := '0';
signal Z28        : std_logic := '0';
signal Z29        : std_logic := '0';
signal Z30        : std_logic := '0';
signal Z31        : std_logic := '0';
signal Z32        : std_logic := '0';
signal Z33        : std_logic := '0';
signal Z34        : std_logic := '0';
signal Z35        : std_logic := '0';
signal Z36        : std_logic := '0';
signal Z37        : std_logic := '0';
signal Z38        : std_logic := '0';
signal Z39        : std_logic := '0';
signal Z40        : std_logic := '0';
signal Z41        : std_logic := '0';
signal Z42        : std_logic := '0';
signal Z43        : std_logic := '0';
signal Z44        : std_logic := '0';
signal Z45        : std_logic := '0';
signal Z46        : std_logic := '0';
signal Z47        : std_logic := '0';
signal Z48        : std_logic := '0';
signal Z49        : std_logic := '0';
signal Z50        : std_logic := '0';
signal Z51        : std_logic := '0';
signal Z52        : std_logic := '0';
signal Z53        : std_logic := '0';
signal Z54        : std_logic := '0';
signal Z55        : std_logic := '0';


constant raw_config0_gen : bit_vector(19 downto 0)
    := CO_SEL & ALU_DYNAMIC_OP & SATURATION_RANK & ENABLE_SATURATION & Z_FEEDBACK_SHL12 & MUX_Z &
       MUX_CI & MUX_Y & MUX_X & MUX_P & MUX_B & MUX_A & PRE_ADDER_OP & SIGNED_MODE;

constant raw_config1_gen : bit_vector(18 downto 0)
    := PR_OV_MUX & PR_CO_MUX & PR_Z_MUX & PR_ALU_MUX & PR_MULT_MUX & PR_Y_MUX & PR_X_MUX &
       PR_P_MUX & PR_CI_MUX & PR_D_MUX & PR_C_MUX & PR_B_CASCADE_MUX & PR_B_MUX & PR_A_CASCADE_MUX &
       PR_A_MUX;

constant raw_config2_gen : bit_vector(12 downto 0)
    := ENABLE_PR_OV_RST & ENABLE_PR_CO_RST & ENABLE_PR_Z_RST & ENABLE_PR_ALU_RST &
       ENABLE_PR_MULT_RST & ENABLE_PR_Y_RST & ENABLE_PR_X_RST & ENABLE_PR_P_RST & ENABLE_PR_CI_RST &
       ENABLE_PR_D_RST & ENABLE_PR_C_RST & ENABLE_PR_B_RST & ENABLE_PR_A_RST;

constant raw_config3_gen : bit_vector(6 downto 0) := ALU_MUX & ALU_OP;


----------------------------------------------------------
-- NX_DSP declaration
----------------------------------------------------------
component NX_DSP
generic (
   std_mode    : string := ""; -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
   raw_config0 : bit_vector(19 downto 0) := B"00000000000000000000";        -- MUX
   raw_config1 : bit_vector(18 downto 0) := B"0000000000000000000";         -- PRC
   raw_config2 : bit_vector(12 downto 0) := B"0000000000000";               -- PRR
   raw_config3 : bit_vector( 6 downto 0) := B"0000000"                      -- ALU
   );
port (
   A1         : in std_logic := '0';
   A2         : in std_logic := '0';
   A3         : in std_logic := '0';
   A4         : in std_logic := '0';
   A5         : in std_logic := '0';
   A6         : in std_logic := '0';
   A7         : in std_logic := '0';
   A8         : in std_logic := '0';
   A9         : in std_logic := '0';
   A10        : in std_logic := '0';
   A11        : in std_logic := '0';
   A12        : in std_logic := '0';
   A13        : in std_logic := '0';
   A14        : in std_logic := '0';
   A15        : in std_logic := '0';
   A16        : in std_logic := '0';
   A17        : in std_logic := '0';
   A18        : in std_logic := '0';
   A19        : in std_logic := '0';
   A20        : in std_logic := '0';
   A21        : in std_logic := '0';
   A22        : in std_logic := '0';
   A23        : in std_logic := '0';
   A24        : in std_logic := '0';

   B1         : in std_logic := '0';
   B2         : in std_logic := '0';
   B3         : in std_logic := '0';
   B4         : in std_logic := '0';
   B5         : in std_logic := '0';
   B6         : in std_logic := '0';
   B7         : in std_logic := '0';
   B8         : in std_logic := '0';
   B9         : in std_logic := '0';
   B10        : in std_logic := '0';
   B11        : in std_logic := '0';
   B12        : in std_logic := '0';
   B13        : in std_logic := '0';
   B14        : in std_logic := '0';
   B15        : in std_logic := '0';
   B16        : in std_logic := '0';
   B17        : in std_logic := '0';
   B18        : in std_logic := '0';

   C1         : in std_logic := '0';
   C2         : in std_logic := '0';
   C3         : in std_logic := '0';
   C4         : in std_logic := '0';
   C5         : in std_logic := '0';
   C6         : in std_logic := '0';
   C7         : in std_logic := '0';
   C8         : in std_logic := '0';
   C9         : in std_logic := '0';
   C10        : in std_logic := '0';
   C11        : in std_logic := '0';
   C12        : in std_logic := '0';
   C13        : in std_logic := '0';
   C14        : in std_logic := '0';
   C15        : in std_logic := '0';
   C16        : in std_logic := '0';
   C17        : in std_logic := '0';
   C18        : in std_logic := '0';
   C19        : in std_logic := '0';
   C20        : in std_logic := '0';
   C21        : in std_logic := '0';
   C22        : in std_logic := '0';
   C23        : in std_logic := '0';
   C24        : in std_logic := '0';
   C25        : in std_logic := '0';
   C26        : in std_logic := '0';
   C27        : in std_logic := '0';
   C28        : in std_logic := '0';
   C29        : in std_logic := '0';
   C30        : in std_logic := '0';
   C31        : in std_logic := '0';
   C32        : in std_logic := '0';
   C33        : in std_logic := '0';
   C34        : in std_logic := '0';
   C35        : in std_logic := '0';
   C36        : in std_logic := '0';

   CAI1       : in std_logic := '0';
   CAI2       : in std_logic := '0';
   CAI3       : in std_logic := '0';
   CAI4       : in std_logic := '0';
   CAI5       : in std_logic := '0';
   CAI6       : in std_logic := '0';
   CAI7       : in std_logic := '0';
   CAI8       : in std_logic := '0';
   CAI9       : in std_logic := '0';
   CAI10      : in std_logic := '0';
   CAI11      : in std_logic := '0';
   CAI12      : in std_logic := '0';
   CAI13      : in std_logic := '0';
   CAI14      : in std_logic := '0';
   CAI15      : in std_logic := '0';
   CAI16      : in std_logic := '0';
   CAI17      : in std_logic := '0';
   CAI18      : in std_logic := '0';

   CAO1       : out std_logic := '0';
   CAO2       : out std_logic := '0';
   CAO3       : out std_logic := '0';
   CAO4       : out std_logic := '0';
   CAO5       : out std_logic := '0';
   CAO6       : out std_logic := '0';
   CAO7       : out std_logic := '0';
   CAO8       : out std_logic := '0';
   CAO9       : out std_logic := '0';
   CAO10      : out std_logic := '0';
   CAO11      : out std_logic := '0';
   CAO12      : out std_logic := '0';
   CAO13      : out std_logic := '0';
   CAO14      : out std_logic := '0';
   CAO15      : out std_logic := '0';
   CAO16      : out std_logic := '0';
   CAO17      : out std_logic := '0';
   CAO18      : out std_logic := '0';

   CBI1       : in std_logic := '0';
   CBI2       : in std_logic := '0';
   CBI3       : in std_logic := '0';
   CBI4       : in std_logic := '0';
   CBI5       : in std_logic := '0';
   CBI6       : in std_logic := '0';
   CBI7       : in std_logic := '0';
   CBI8       : in std_logic := '0';
   CBI9       : in std_logic := '0';
   CBI10      : in std_logic := '0';
   CBI11      : in std_logic := '0';
   CBI12      : in std_logic := '0';
   CBI13      : in std_logic := '0';
   CBI14      : in std_logic := '0';
   CBI15      : in std_logic := '0';
   CBI16      : in std_logic := '0';
   CBI17      : in std_logic := '0';
   CBI18      : in std_logic := '0';

   CBO1       : out std_logic := '0';
   CBO2       : out std_logic := '0';
   CBO3       : out std_logic := '0';
   CBO4       : out std_logic := '0';
   CBO5       : out std_logic := '0';
   CBO6       : out std_logic := '0';
   CBO7       : out std_logic := '0';
   CBO8       : out std_logic := '0';
   CBO9       : out std_logic := '0';
   CBO10      : out std_logic := '0';
   CBO11      : out std_logic := '0';
   CBO12      : out std_logic := '0';
   CBO13      : out std_logic := '0';
   CBO14      : out std_logic := '0';
   CBO15      : out std_logic := '0';
   CBO16      : out std_logic := '0';
   CBO17      : out std_logic := '0';
   CBO18      : out std_logic := '0';

   CCI        : in std_logic := '0';
   CCO        : out std_logic := '0';
   CI         : in std_logic := '0';
   CK         : in std_logic := '0';
   CO         : out std_logic := '0';
   CO37       : out std_logic := '0';
   CO49       : out std_logic := '0';

   CZI1       : in std_logic := '0';
   CZI2       : in std_logic := '0';
   CZI3       : in std_logic := '0';
   CZI4       : in std_logic := '0';
   CZI5       : in std_logic := '0';
   CZI6       : in std_logic := '0';
   CZI7       : in std_logic := '0';
   CZI8       : in std_logic := '0';
   CZI9       : in std_logic := '0';
   CZI10      : in std_logic := '0';
   CZI11      : in std_logic := '0';
   CZI12      : in std_logic := '0';
   CZI13      : in std_logic := '0';
   CZI14      : in std_logic := '0';
   CZI15      : in std_logic := '0';
   CZI16      : in std_logic := '0';
   CZI17      : in std_logic := '0';
   CZI18      : in std_logic := '0';
   CZI19      : in std_logic := '0';
   CZI20      : in std_logic := '0';
   CZI21      : in std_logic := '0';
   CZI22      : in std_logic := '0';
   CZI23      : in std_logic := '0';
   CZI24      : in std_logic := '0';
   CZI25      : in std_logic := '0';
   CZI26      : in std_logic := '0';
   CZI27      : in std_logic := '0';
   CZI28      : in std_logic := '0';
   CZI29      : in std_logic := '0';
   CZI30      : in std_logic := '0';
   CZI31      : in std_logic := '0';
   CZI32      : in std_logic := '0';
   CZI33      : in std_logic := '0';
   CZI34      : in std_logic := '0';
   CZI35      : in std_logic := '0';
   CZI36      : in std_logic := '0';
   CZI37      : in std_logic := '0';
   CZI38      : in std_logic := '0';
   CZI39      : in std_logic := '0';
   CZI40      : in std_logic := '0';
   CZI41      : in std_logic := '0';
   CZI42      : in std_logic := '0';
   CZI43      : in std_logic := '0';
   CZI44      : in std_logic := '0';
   CZI45      : in std_logic := '0';
   CZI46      : in std_logic := '0';
   CZI47      : in std_logic := '0';
   CZI48      : in std_logic := '0';
   CZI49      : in std_logic := '0';
   CZI50      : in std_logic := '0';
   CZI51      : in std_logic := '0';
   CZI52      : in std_logic := '0';
   CZI53      : in std_logic := '0';
   CZI54      : in std_logic := '0';
   CZI55      : in std_logic := '0';
   CZI56      : in std_logic := '0';

   CZO1       : out std_logic := '0';
   CZO2       : out std_logic := '0';
   CZO3       : out std_logic := '0';
   CZO4       : out std_logic := '0';
   CZO5       : out std_logic := '0';
   CZO6       : out std_logic := '0';
   CZO7       : out std_logic := '0';
   CZO8       : out std_logic := '0';
   CZO9       : out std_logic := '0';
   CZO10      : out std_logic := '0';
   CZO11      : out std_logic := '0';
   CZO12      : out std_logic := '0';
   CZO13      : out std_logic := '0';
   CZO14      : out std_logic := '0';
   CZO15      : out std_logic := '0';
   CZO16      : out std_logic := '0';
   CZO17      : out std_logic := '0';
   CZO18      : out std_logic := '0';
   CZO19      : out std_logic := '0';
   CZO20      : out std_logic := '0';
   CZO21      : out std_logic := '0';
   CZO22      : out std_logic := '0';
   CZO23      : out std_logic := '0';
   CZO24      : out std_logic := '0';
   CZO25      : out std_logic := '0';
   CZO26      : out std_logic := '0';
   CZO27      : out std_logic := '0';
   CZO28      : out std_logic := '0';
   CZO29      : out std_logic := '0';
   CZO30      : out std_logic := '0';
   CZO31      : out std_logic := '0';
   CZO32      : out std_logic := '0';
   CZO33      : out std_logic := '0';
   CZO34      : out std_logic := '0';
   CZO35      : out std_logic := '0';
   CZO36      : out std_logic := '0';
   CZO37      : out std_logic := '0';
   CZO38      : out std_logic := '0';
   CZO39      : out std_logic := '0';
   CZO40      : out std_logic := '0';
   CZO41      : out std_logic := '0';
   CZO42      : out std_logic := '0';
   CZO43      : out std_logic := '0';
   CZO44      : out std_logic := '0';
   CZO45      : out std_logic := '0';
   CZO46      : out std_logic := '0';
   CZO47      : out std_logic := '0';
   CZO48      : out std_logic := '0';
   CZO49      : out std_logic := '0';
   CZO50      : out std_logic := '0';
   CZO51      : out std_logic := '0';
   CZO52      : out std_logic := '0';
   CZO53      : out std_logic := '0';
   CZO54      : out std_logic := '0';
   CZO55      : out std_logic := '0';
   CZO56      : out std_logic := '0';

   D1         : in std_logic := '0';
   D2         : in std_logic := '0';
   D3         : in std_logic := '0';
   D4         : in std_logic := '0';
   D5         : in std_logic := '0';
   D6         : in std_logic := '0';
   D7         : in std_logic := '0';
   D8         : in std_logic := '0';
   D9         : in std_logic := '0';
   D10        : in std_logic := '0';
   D11        : in std_logic := '0';
   D12        : in std_logic := '0';
   D13        : in std_logic := '0';
   D14        : in std_logic := '0';
   D15        : in std_logic := '0';
   D16        : in std_logic := '0';
   D17        : in std_logic := '0';
   D18        : in std_logic := '0';

   OVF        : out std_logic := '0';
   R          : in std_logic := '0';
   RZ         : in std_logic := '0';
   WE         : in std_logic := '0';

   Z1         : out std_logic := '0';
   Z2         : out std_logic := '0';
   Z3         : out std_logic := '0';
   Z4         : out std_logic := '0';
   Z5         : out std_logic := '0';
   Z6         : out std_logic := '0';
   Z7         : out std_logic := '0';
   Z8         : out std_logic := '0';
   Z9         : out std_logic := '0';
   Z10        : out std_logic := '0';
   Z11        : out std_logic := '0';
   Z12        : out std_logic := '0';
   Z13        : out std_logic := '0';
   Z14        : out std_logic := '0';
   Z15        : out std_logic := '0';
   Z16        : out std_logic := '0';
   Z17        : out std_logic := '0';
   Z18        : out std_logic := '0';
   Z19        : out std_logic := '0';
   Z20        : out std_logic := '0';
   Z21        : out std_logic := '0';
   Z22        : out std_logic := '0';
   Z23        : out std_logic := '0';
   Z24        : out std_logic := '0';
   Z25        : out std_logic := '0';
   Z26        : out std_logic := '0';
   Z27        : out std_logic := '0';
   Z28        : out std_logic := '0';
   Z29        : out std_logic := '0';
   Z30        : out std_logic := '0';
   Z31        : out std_logic := '0';
   Z32        : out std_logic := '0';
   Z33        : out std_logic := '0';
   Z34        : out std_logic := '0';
   Z35        : out std_logic := '0';
   Z36        : out std_logic := '0';
   Z37        : out std_logic := '0';
   Z38        : out std_logic := '0';
   Z39        : out std_logic := '0';
   Z40        : out std_logic := '0';
   Z41        : out std_logic := '0';
   Z42        : out std_logic := '0';
   Z43        : out std_logic := '0';
   Z44        : out std_logic := '0';
   Z45        : out std_logic := '0';
   Z46        : out std_logic := '0';
   Z47        : out std_logic := '0';
   Z48        : out std_logic := '0';
   Z49        : out std_logic := '0';
   Z50        : out std_logic := '0';
   Z51        : out std_logic := '0';
   Z52        : out std_logic := '0';
   Z53        : out std_logic := '0';
   Z54        : out std_logic := '0';
   Z55        : out std_logic := '0';
   Z56        : out std_logic := '0'
   );
end component;

begin

----------------------------------------------------------
-- Instantiation the NX_DSP component
----------------------------------------------------------
DSP_INST : NX_DSP
generic map (
   std_mode    => "", -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
   raw_config0 => raw_config0_gen, -- MODE and MUXes
   raw_config1 => raw_config1_gen, -- Pipeline Registers
   raw_config2 => raw_config2_gen, -- Reset Enable for internal registers
   raw_config3 => raw_config3_gen   -- ALU modes
   )
port map (
   A1         => A(0),
   A2         => A(1),
   A3         => A(2),
   A4         => A(3),
   A5         => A(4),
   A6         => A(5),
   A7         => A(6),
   A8         => A(7),
   A9         => A(8),
   A10        => A(9),
   A11        => A(10),
   A12        => A(11),
   A13        => A(12),
   A14        => A(13),
   A15        => A(14),
   A16        => A(15),
   A17        => A(16),
   A18        => A(17),
   A19        => A(18),
   A20        => A(19),
   A21        => A(20),
   A22        => A(21),
   A23        => A(22),
   A24        => A(23),

   B1         => B(0),
   B2         => B(1),
   B3         => B(2),
   B4         => B(3),
   B5         => B(4),
   B6         => B(5),
   B7         => B(6),
   B8         => B(7),
   B9         => B(8),
   B10        => B(9),
   B11        => B(10),
   B12        => B(11),
   B13        => B(12),
   B14        => B(13),
   B15        => B(14),
   B16        => B(15),
   B17        => B(16),
   B18        => B(17),

   C1         => C(0),
   C2         => C(1),
   C3         => C(2),
   C4         => C(3),
   C5         => C(4),
   C6         => C(5),
   C7         => C(6),
   C8         => C(7),
   C9         => C(8),
   C10        => C(9),
   C11        => C(10),
   C12        => C(11),
   C13        => C(12),
   C14        => C(13),
   C15        => C(14),
   C16        => C(15),
   C17        => C(16),
   C18        => C(17),
   C19        => C(18),
   C20        => C(19),
   C21        => C(20),
   C22        => C(21),
   C23        => C(22),
   C24        => C(23),
   C25        => C(24),
   C26        => C(25),
   C27        => C(26),
   C28        => C(27),
   C29        => C(28),
   C30        => C(29),
   C31        => C(30),
   C32        => C(31),
   C33        => C(32),
   C34        => C(33),
   C35        => C(34),
   C36        => C(35),

   CAI1       => CAI(0),
   CAI2       => CAI(1),
   CAI3       => CAI(2),
   CAI4       => CAI(3),
   CAI5       => CAI(4),
   CAI6       => CAI(5),
   CAI7       => CAI(6),
   CAI8       => CAI(7),
   CAI9       => CAI(8),
   CAI10      => CAI(9),
   CAI11      => CAI(10),
   CAI12      => CAI(11),
   CAI13      => CAI(12),
   CAI14      => CAI(13),
   CAI15      => CAI(14),
   CAI16      => CAI(15),
   CAI17      => CAI(16),
   CAI18      => CAI(17),

   CAO1       => CAO(0),
   CAO2       => CAO(1),
   CAO3       => CAO(2),
   CAO4       => CAO(3),
   CAO5       => CAO(4),
   CAO6       => CAO(5),
   CAO7       => CAO(6),
   CAO8       => CAO(7),
   CAO9       => CAO(8),
   CAO10      => CAO(9),
   CAO11      => CAO(10),
   CAO12      => CAO(11),
   CAO13      => CAO(12),
   CAO14      => CAO(13),
   CAO15      => CAO(14),
   CAO16      => CAO(15),
   CAO17      => CAO(16),
   CAO18      => CAO(17),

   CBI1       => CBI(0),
   CBI2       => CBI(1),
   CBI3       => CBI(2),
   CBI4       => CBI(3),
   CBI5       => CBI(4),
   CBI6       => CBI(5),
   CBI7       => CBI(6),
   CBI8       => CBI(7),
   CBI9       => CBI(8),
   CBI10      => CBI(9),
   CBI11      => CBI(10),
   CBI12      => CBI(11),
   CBI13      => CBI(12),
   CBI14      => CBI(13),
   CBI15      => CBI(14),
   CBI16      => CBI(15),
   CBI17      => CBI(16),
   CBI18      => CBI(17),

   CBO1       => CBO(0),
   CBO2       => CBO(1),
   CBO3       => CBO(2),
   CBO4       => CBO(3),
   CBO5       => CBO(4),
   CBO6       => CBO(5),
   CBO7       => CBO(6),
   CBO8       => CBO(7),
   CBO9       => CBO(8),
   CBO10      => CBO(9),
   CBO11      => CBO(10),
   CBO12      => CBO(11),
   CBO13      => CBO(12),
   CBO14      => CBO(13),
   CBO15      => CBO(14),
   CBO16      => CBO(15),
   CBO17      => CBO(16),
   CBO18      => CBO(17),

   CCI        => CCI,
   CCO        => CCO,
   CI         => CI,
   CK         => CK,
   CO         => CO,
   CO37       => CO36,
   CO49       => CO48,

   CZI1       => CZI(0),
   CZI2       => CZI(1),
   CZI3       => CZI(2),
   CZI4       => CZI(3),
   CZI5       => CZI(4),
   CZI6       => CZI(5),
   CZI7       => CZI(6),
   CZI8       => CZI(7),
   CZI9       => CZI(8),
   CZI10      => CZI(9),
   CZI11      => CZI(10),
   CZI12      => CZI(11),
   CZI13      => CZI(12),
   CZI14      => CZI(13),
   CZI15      => CZI(14),
   CZI16      => CZI(15),
   CZI17      => CZI(16),
   CZI18      => CZI(17),
   CZI19      => CZI(18),
   CZI20      => CZI(19),
   CZI21      => CZI(20),
   CZI22      => CZI(21),
   CZI23      => CZI(22),
   CZI24      => CZI(23),
   CZI25      => CZI(24),
   CZI26      => CZI(25),
   CZI27      => CZI(26),
   CZI28      => CZI(27),
   CZI29      => CZI(28),
   CZI30      => CZI(29),
   CZI31      => CZI(30),
   CZI32      => CZI(31),
   CZI33      => CZI(32),
   CZI34      => CZI(33),
   CZI35      => CZI(34),
   CZI36      => CZI(35),
   CZI37      => CZI(36),
   CZI38      => CZI(37),
   CZI39      => CZI(38),
   CZI40      => CZI(39),
   CZI41      => CZI(40),
   CZI42      => CZI(41),
   CZI43      => CZI(42),
   CZI44      => CZI(43),
   CZI45      => CZI(44),
   CZI46      => CZI(45),
   CZI47      => CZI(46),
   CZI48      => CZI(47),
   CZI49      => CZI(48),
   CZI50      => CZI(49),
   CZI51      => CZI(50),
   CZI52      => CZI(51),
   CZI53      => CZI(52),
   CZI54      => CZI(53),
   CZI55      => CZI(54),
   CZI56      => CZI(55),

   CZO1       => CZO(0),
   CZO2       => CZO(1),
   CZO3       => CZO(2),
   CZO4       => CZO(3),
   CZO5       => CZO(4),
   CZO6       => CZO(5),
   CZO7       => CZO(6),
   CZO8       => CZO(7),
   CZO9       => CZO(8),
   CZO10      => CZO(9),
   CZO11      => CZO(10),
   CZO12      => CZO(11),
   CZO13      => CZO(12),
   CZO14      => CZO(13),
   CZO15      => CZO(14),
   CZO16      => CZO(15),
   CZO17      => CZO(16),
   CZO18      => CZO(17),
   CZO19      => CZO(18),
   CZO20      => CZO(19),
   CZO21      => CZO(20),
   CZO22      => CZO(21),
   CZO23      => CZO(22),
   CZO24      => CZO(23),
   CZO25      => CZO(24),
   CZO26      => CZO(25),
   CZO27      => CZO(26),
   CZO28      => CZO(27),
   CZO29      => CZO(28),
   CZO30      => CZO(29),
   CZO31      => CZO(30),
   CZO32      => CZO(31),
   CZO33      => CZO(32),
   CZO34      => CZO(33),
   CZO35      => CZO(34),
   CZO36      => CZO(35),
   CZO37      => CZO(36),
   CZO38      => CZO(37),
   CZO39      => CZO(38),
   CZO40      => CZO(39),
   CZO41      => CZO(40),
   CZO42      => CZO(41),
   CZO43      => CZO(42),
   CZO44      => CZO(43),
   CZO45      => CZO(44),
   CZO46      => CZO(45),
   CZO47      => CZO(46),
   CZO48      => CZO(47),
   CZO49      => CZO(48),
   CZO50      => CZO(49),
   CZO51      => CZO(50),
   CZO52      => CZO(51),
   CZO53      => CZO(52),
   CZO54      => CZO(53),
   CZO55      => CZO(54),
   CZO56      => CZO(55),

   D1         => D(0),
   D2         => D(1),
   D3         => D(2),
   D4         => D(3),
   D5         => D(4),
   D6         => D(5),
   D7         => D(6),
   D8         => D(7),
   D9         => D(8),
   D10        => D(9),
   D11        => D(10),
   D12        => D(11),
   D13        => D(12),
   D14        => D(13),
   D15        => D(14),
   D16        => D(15),
   D17        => D(16),
   D18        => D(17),

   OVF        => OVF,
   R          => R,
   RZ         => RZ,
   WE         => WE,

   Z1         => Z(0),
   Z2         => Z(1),
   Z3         => Z(2),
   Z4         => Z(3),
   Z5         => Z(4),
   Z6         => Z(5),
   Z7         => Z(6),
   Z8         => Z(7),
   Z9         => Z(8),
   Z10        => Z(9),
   Z11        => Z(10),
   Z12        => Z(11),
   Z13        => Z(12),
   Z14        => Z(13),
   Z15        => Z(14),
   Z16        => Z(15),
   Z17        => Z(16),
   Z18        => Z(17),
   Z19        => Z(18),
   Z20        => Z(19),
   Z21        => Z(20),
   Z22        => Z(21),
   Z23        => Z(22),
   Z24        => Z(23),
   Z25        => Z(24),
   Z26        => Z(25),
   Z27        => Z(26),
   Z28        => Z(27),
   Z29        => Z(28),
   Z30        => Z(29),
   Z31        => Z(30),
   Z32        => Z(31),
   Z33        => Z(32),
   Z34        => Z(33),
   Z35        => Z(34),
   Z36        => Z(35),
   Z37        => Z(36),
   Z38        => Z(37),
   Z39        => Z(38),
   Z40        => Z(39),
   Z41        => Z(40),
   Z42        => Z(41),
   Z43        => Z(42),
   Z44        => Z(43),
   Z45        => Z(44),
   Z46        => Z(45),
   Z47        => Z(46),
   Z48        => Z(47),
   Z49        => Z(48),
   Z50        => Z(49),
   Z51        => Z(50),
   Z52        => Z(51),
   Z53        => Z(52),
   Z54        => Z(53),
   Z55        => Z(54),
   Z56        => Z(55)
   );

end NX_RTL;
-- #}}}#
-- =================================================================================================
--   NX_DSPDPRAM_FULL_U definition                                                       2020/02/03
-- =================================================================================================

-- NX_DSPDPRAM_FULL_U#{{{#
library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DSPDPRAM_FULL_U is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    dsp0_clk_i  : in  std_logic;                                        -- DSP1.CK
    dsp0_rst_i  : in  std_logic; -- rst_i  et rstsys_i                  -- DSP1.R
    dsp0_rstz_i : in  std_logic; -- rstz_i et rstzsys_i                 -- DSP1.RZ
    dsp0_we_i   : in  std_logic; -- we_i   et wesys_i                   -- DSP1.WE
    dsp0_wez_i  : in  std_logic; -- wez_i  et wezsys_i                  -- DSP1.WEZ
    dsp0_cy_i   : in  std_logic;                                        -- DSP1.CI
    dsp0_a_i    : in  std_logic_vector(23 downto 0);                    -- DSP1.A
    dsp0_b_i    : in  std_logic_vector(17 downto 0);                    -- DSP1.B
    dsp0_c_i    : in  std_logic_vector(35 downto 0);                    -- DSP1.C
    dsp0_d_i    : in  std_logic_vector(17 downto 0);                    -- DSP1.D

    dsp0_z_o    : out std_logic_vector(55 downto 0);                    -- DSP1.Z
    dsp0_cy_o   : out std_logic;                                        -- DSP1.RESERVED
    dsp0_cy42_o : out std_logic;                                        -- DSP1.CO43
    dsp0_cy56_o : out std_logic;                                        -- DSP1.CO57
    dsp0_ovf_o  : out std_logic;                                        -- DSP1.OVF

    dsp1_clk_i  : in  std_logic;                                        -- DSP2.CK
    dsp1_rst_i  : in  std_logic; -- rst_i  et rstsys_i                  -- DSP2.R
    dsp1_rstz_i : in  std_logic; -- rstz_i et rstzsys_i                 -- DSP2.RZ
    dsp1_we_i   : in  std_logic; -- we_i   et wesys_i                   -- DSP2.WE
    dsp1_wez_i  : in  std_logic; -- wez_i  et wezsys_i                  -- DSP2.WE
    dsp1_cy_i   : in  std_logic;                                        -- DSP2.CI
    dsp1_a_i    : in  std_logic_vector(23 downto 0);                    -- DSP2.A
    dsp1_b_i    : in  std_logic_vector(17 downto 0);                    -- DSP2.B
    dsp1_c_i    : in  std_logic_vector(35 downto 0);                    -- DSP2.C
    dsp1_d_i    : in  std_logic_vector(17 downto 0);                    -- DSP2.D

    dsp1_z_o    : out std_logic_vector(55 downto 0);                    -- DSP2.Z
    dsp1_cy_o   : out std_logic;                                        -- DSP2.RESERVED
    dsp1_cy42_o : out std_logic;                                        -- DSP2.CO43
    dsp1_cy56_o : out std_logic;                                        -- DSP2.CO57
    dsp1_ovf_o  : out std_logic;                                        -- DSP2.OVF

    dpram_clkmem0_i          : in  std_logic;                           -- RAM.ACK
    dpram_rst0_i             : in  std_logic; -- rst_i et rstsys_i      -- RAM.AR
    dpram_cs0_i              : in  std_logic; -- cs_i  et cssys_i       -- RAM.ACS
    dpram_we0_i              : in  std_logic; -- we_i  et wesys_i       -- RAM.AWE
    dpram_addr0_i            : in  std_logic_vector(15 downto 0);       -- RAM.AA
    dpram_din0_i             : in  std_logic_vector(23 downto 0);       -- RAM.AI
    dpram_dout0_o            : out std_logic_vector(23 downto 0);       -- RAM.AO
    dpram_ecc_corrected0_o   : out std_logic;                           -- RAM.ACOR
    dpram_ecc_uncorrected0_o : out std_logic;                           -- RAM.AERR

    dpram_clkmem1_i          : in  std_logic;                           -- RAM.BCK
    dpram_rst1_i             : in  std_logic; -- rst_i et rstsys_i      -- RAM.BR
    dpram_cs1_i              : in  std_logic; -- cs_i  et cssys_i       -- RAM.BCS
    dpram_we1_i              : in  std_logic; -- we_i  et wesys_i       -- RAM.BWE
    dpram_addr1_i            : in  std_logic_vector(15 downto 0);       -- RAM.BA
    dpram_din1_i             : in  std_logic_vector(23 downto 0);       -- RAM.BI
    dpram_dout1_o            : out std_logic_vector(23 downto 0);       -- RAM.BO
    dpram_ecc_corrected1_o   : out std_logic;                           -- RAM.BCOR
    dpram_ecc_uncorrected1_o : out std_logic                            -- RAM.BERR
);
end NX_DSPDPRAM_FULL_U;
--#}}}#

-- architecture NX_RTL of NX_DSPDPRAM_FULL_U#{{{#
architecture NX_RTL of NX_DSPDPRAM_FULL_U is

  -- component NX_DSP_U_BOX#{{{#
  component NX_DSP_U_BOX
  generic (
      col    : integer := 2;
      row    : integer := 6;
      cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
      cfg_top_i : bit_vector(95 downto 0) := (others => '0')
  );
  port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    RESERVED: out std_logic;
    CO43  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;
    WEZ   : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
  );
  end component;
  --#}}}#

  -- component NX_RAM_U_BOX#{{{#
  component NX_RAM_U_BOX
  generic (
      col    : integer := 2;
      row    : integer := 6;
      cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
      cfg_top_i : bit_vector(95 downto 0) := (others => '0')
  );
  port (
    ACK   : in  std_logic;
    BCK   : in  std_logic;

    AI1   : in  std_logic;
    AI2   : in  std_logic;
    AI3   : in  std_logic;
    AI4   : in  std_logic;
    AI5   : in  std_logic;
    AI6   : in  std_logic;
    AI7   : in  std_logic;
    AI8   : in  std_logic;
    AI9   : in  std_logic;
    AI10  : in  std_logic;
    AI11  : in  std_logic;
    AI12  : in  std_logic;
    AI13  : in  std_logic;
    AI14  : in  std_logic;
    AI15  : in  std_logic;
    AI16  : in  std_logic;
    AI17  : in  std_logic;
    AI18  : in  std_logic;
    AI19  : in  std_logic;
    AI20  : in  std_logic;
    AI21  : in  std_logic;
    AI22  : in  std_logic;
    AI23  : in  std_logic;
    AI24  : in  std_logic;

    BI1   : in  std_logic;
    BI2   : in  std_logic;
    BI3   : in  std_logic;
    BI4   : in  std_logic;
    BI5   : in  std_logic;
    BI6   : in  std_logic;
    BI7   : in  std_logic;
    BI8   : in  std_logic;
    BI9   : in  std_logic;
    BI10  : in  std_logic;
    BI11  : in  std_logic;
    BI12  : in  std_logic;
    BI13  : in  std_logic;
    BI14  : in  std_logic;
    BI15  : in  std_logic;
    BI16  : in  std_logic;
    BI17  : in  std_logic;
    BI18  : in  std_logic;
    BI19  : in  std_logic;
    BI20  : in  std_logic;
    BI21  : in  std_logic;
    BI22  : in  std_logic;
    BI23  : in  std_logic;
    BI24  : in  std_logic;

    ACOR  : out std_logic;
    AERR  : out std_logic;
    BCOR  : out std_logic;
    BERR  : out std_logic;

    AO1   : out std_logic;
    AO2   : out std_logic;
    AO3   : out std_logic;
    AO4   : out std_logic;
    AO5   : out std_logic;
    AO6   : out std_logic;
    AO7   : out std_logic;
    AO8   : out std_logic;
    AO9   : out std_logic;
    AO10  : out std_logic;
    AO11  : out std_logic;
    AO12  : out std_logic;
    AO13  : out std_logic;
    AO14  : out std_logic;
    AO15  : out std_logic;
    AO16  : out std_logic;
    AO17  : out std_logic;
    AO18  : out std_logic;
    AO19  : out std_logic;
    AO20  : out std_logic;
    AO21  : out std_logic;
    AO22  : out std_logic;
    AO23  : out std_logic;
    AO24  : out std_logic;

    BO1   : out std_logic;
    BO2   : out std_logic;
    BO3   : out std_logic;
    BO4   : out std_logic;
    BO5   : out std_logic;
    BO6   : out std_logic;
    BO7   : out std_logic;
    BO8   : out std_logic;
    BO9   : out std_logic;
    BO10  : out std_logic;
    BO11  : out std_logic;
    BO12  : out std_logic;
    BO13  : out std_logic;
    BO14  : out std_logic;
    BO15  : out std_logic;
    BO16  : out std_logic;
    BO17  : out std_logic;
    BO18  : out std_logic;
    BO19  : out std_logic;
    BO20  : out std_logic;
    BO21  : out std_logic;
    BO22  : out std_logic;
    BO23  : out std_logic;
    BO24  : out std_logic;

    AA1   : in  std_logic;
    AA2   : in  std_logic;
    AA3   : in  std_logic;
    AA4   : in  std_logic;
    AA5   : in  std_logic;
    AA6   : in  std_logic;
    AA7   : in  std_logic;
    AA8   : in  std_logic;
    AA9   : in  std_logic;
    AA10  : in  std_logic;
    AA11  : in  std_logic;
    AA12  : in  std_logic;
    AA13  : in  std_logic;
    AA14  : in  std_logic;
    AA15  : in  std_logic;
    AA16  : in  std_logic;

    ACS   : in  std_logic;
    AWE   : in  std_logic;
    AR    : in  std_logic;

    BA1   : in  std_logic;
    BA2   : in  std_logic;
    BA3   : in  std_logic;
    BA4   : in  std_logic;
    BA5   : in  std_logic;
    BA6   : in  std_logic;
    BA7   : in  std_logic;
    BA8   : in  std_logic;
    BA9   : in  std_logic;
    BA10  : in  std_logic;
    BA11  : in  std_logic;
    BA12  : in  std_logic;
    BA13  : in  std_logic;
    BA14  : in  std_logic;
    BA15  : in  std_logic;
    BA16  : in  std_logic;

    BCS   : in  std_logic;
    BWE   : in  std_logic;
    BR    : in  std_logic
  );
  end component;
  --#}}}#

signal c_cy_int : std_logic;
signal c_a_int : std_logic_vector(23 downto 0);
signal c_b_int : std_logic_vector(17 downto 0);
signal c_z_int : std_logic_vector(55 downto 0);

attribute syn_preserve : boolean;
attribute syn_preserve of dsp_0 : label is true;
attribute syn_preserve of dsp_1 : label is true;
attribute syn_preserve of ram_0 : label is true;

begin

-- instance dsp0#{{{#
dsp_0 : NX_DSP_U_BOX
generic map (
    col    => col
  , row    => row
  , cfg_bot_i => cfg_bot_i
  , cfg_top_i => cfg_top_i
)
port map (
      A1    => dsp0_a_i(0)
   ,  A2    => dsp0_a_i(1)
   ,  A3    => dsp0_a_i(2)
   ,  A4    => dsp0_a_i(3)
   ,  A5    => dsp0_a_i(4)
   ,  A6    => dsp0_a_i(5)
   ,  A7    => dsp0_a_i(6)
   ,  A8    => dsp0_a_i(7)
   ,  A9    => dsp0_a_i(8)
   ,  A10   => dsp0_a_i(9)
   ,  A11   => dsp0_a_i(10)
   ,  A12   => dsp0_a_i(11)
   ,  A13   => dsp0_a_i(12)
   ,  A14   => dsp0_a_i(13)
   ,  A15   => dsp0_a_i(14)
   ,  A16   => dsp0_a_i(15)
   ,  A17   => dsp0_a_i(16)
   ,  A18   => dsp0_a_i(17)
   ,  A19   => dsp0_a_i(18)
   ,  A20   => dsp0_a_i(19)
   ,  A21   => dsp0_a_i(20)
   ,  A22   => dsp0_a_i(21)
   ,  A23   => dsp0_a_i(22)
   ,  A24   => dsp0_a_i(23)
   ,  B1    => dsp0_b_i(0)
   ,  B2    => dsp0_b_i(1)
   ,  B3    => dsp0_b_i(2)
   ,  B4    => dsp0_b_i(3)
   ,  B5    => dsp0_b_i(4)
   ,  B6    => dsp0_b_i(5)
   ,  B7    => dsp0_b_i(6)
   ,  B8    => dsp0_b_i(7)
   ,  B9    => dsp0_b_i(8)
   ,  B10   => dsp0_b_i(9)
   ,  B11   => dsp0_b_i(10)
   ,  B12   => dsp0_b_i(11)
   ,  B13   => dsp0_b_i(12)
   ,  B14   => dsp0_b_i(13)
   ,  B15   => dsp0_b_i(14)
   ,  B16   => dsp0_b_i(15)
   ,  B17   => dsp0_b_i(16)
   ,  B18   => dsp0_b_i(17)
   ,  C1    => dsp0_c_i(0)
   ,  C2    => dsp0_c_i(1)
   ,  C3    => dsp0_c_i(2)
   ,  C4    => dsp0_c_i(3)
   ,  C5    => dsp0_c_i(4)
   ,  C6    => dsp0_c_i(5)
   ,  C7    => dsp0_c_i(6)
   ,  C8    => dsp0_c_i(7)
   ,  C9    => dsp0_c_i(8)
   ,  C10   => dsp0_c_i(9)
   ,  C11   => dsp0_c_i(10)
   ,  C12   => dsp0_c_i(11)
   ,  C13   => dsp0_c_i(12)
   ,  C14   => dsp0_c_i(13)
   ,  C15   => dsp0_c_i(14)
   ,  C16   => dsp0_c_i(15)
   ,  C17   => dsp0_c_i(16)
   ,  C18   => dsp0_c_i(17)
   ,  C19   => dsp0_c_i(18)
   ,  C20   => dsp0_c_i(19)
   ,  C21   => dsp0_c_i(20)
   ,  C22   => dsp0_c_i(21)
   ,  C23   => dsp0_c_i(22)
   ,  C24   => dsp0_c_i(23)
   ,  C25   => dsp0_c_i(24)
   ,  C26   => dsp0_c_i(25)
   ,  C27   => dsp0_c_i(26)
   ,  C28   => dsp0_c_i(27)
   ,  C29   => dsp0_c_i(28)
   ,  C30   => dsp0_c_i(29)
   ,  C31   => dsp0_c_i(30)
   ,  C32   => dsp0_c_i(31)
   ,  C33   => dsp0_c_i(32)
   ,  C34   => dsp0_c_i(33)
   ,  C35   => dsp0_c_i(34)
   ,  C36   => dsp0_c_i(35)
   ,  CAI1  => c_a_int(0)
   ,  CAI2  => c_a_int(1)
   ,  CAI3  => c_a_int(2)
   ,  CAI4  => c_a_int(3)
   ,  CAI5  => c_a_int(4)
   ,  CAI6  => c_a_int(5)
   ,  CAI7  => c_a_int(6)
   ,  CAI8  => c_a_int(7)
   ,  CAI9  => c_a_int(8)
   ,  CAI10 => c_a_int(9)
   ,  CAI11 => c_a_int(10)
   ,  CAI12 => c_a_int(11)
   ,  CAI13 => c_a_int(12)
   ,  CAI14 => c_a_int(13)
   ,  CAI15 => c_a_int(14)
   ,  CAI16 => c_a_int(15)
   ,  CAI17 => c_a_int(16)
   ,  CAI18 => c_a_int(17)
   ,  CAI19 => c_a_int(18)
   ,  CAI20 => c_a_int(19)
   ,  CAI21 => c_a_int(20)
   ,  CAI22 => c_a_int(21)
   ,  CAI23 => c_a_int(22)
   ,  CAI24 => c_a_int(23)
   ,  CAO1  => OPEN
   ,  CAO2  => OPEN
   ,  CAO3  => OPEN
   ,  CAO4  => OPEN
   ,  CAO5  => OPEN
   ,  CAO6  => OPEN
   ,  CAO7  => OPEN
   ,  CAO8  => OPEN
   ,  CAO9  => OPEN
   ,  CAO10 => OPEN
   ,  CAO11 => OPEN
   ,  CAO12 => OPEN
   ,  CAO13 => OPEN
   ,  CAO14 => OPEN
   ,  CAO15 => OPEN
   ,  CAO16 => OPEN
   ,  CAO17 => OPEN
   ,  CAO18 => OPEN
   ,  CAO19 => OPEN
   ,  CAO20 => OPEN
   ,  CAO21 => OPEN
   ,  CAO22 => OPEN
   ,  CAO23 => OPEN
   ,  CAO24 => OPEN
   ,  CBI1  => c_b_int(0)
   ,  CBI2  => c_b_int(1)
   ,  CBI3  => c_b_int(2)
   ,  CBI4  => c_b_int(3)
   ,  CBI5  => c_b_int(4)
   ,  CBI6  => c_b_int(5)
   ,  CBI7  => c_b_int(6)
   ,  CBI8  => c_b_int(7)
   ,  CBI9  => c_b_int(8)
   ,  CBI10 => c_b_int(9)
   ,  CBI11 => c_b_int(10)
   ,  CBI12 => c_b_int(11)
   ,  CBI13 => c_b_int(12)
   ,  CBI14 => c_b_int(13)
   ,  CBI15 => c_b_int(14)
   ,  CBI16 => c_b_int(15)
   ,  CBI17 => c_b_int(16)
   ,  CBI18 => c_b_int(17)
   ,  CBO1  => OPEN
   ,  CBO2  => OPEN
   ,  CBO3  => OPEN
   ,  CBO4  => OPEN
   ,  CBO5  => OPEN
   ,  CBO6  => OPEN
   ,  CBO7  => OPEN
   ,  CBO8  => OPEN
   ,  CBO9  => OPEN
   ,  CBO10 => OPEN
   ,  CBO11 => OPEN
   ,  CBO12 => OPEN
   ,  CBO13 => OPEN
   ,  CBO14 => OPEN
   ,  CBO15 => OPEN
   ,  CBO16 => OPEN
   ,  CBO17 => OPEN
   ,  CBO18 => OPEN
   ,  CCI   => '0'
   ,  CCO   => c_cy_int
   ,  CI    => dsp0_cy_i
   ,  CK    => dsp0_clk_i
   ,  RESERVED => dsp0_cy_o
   ,  CO43  => dsp0_cy42_o
   ,  CO57  => dsp0_cy56_o
   ,  CZI1  => c_z_int(0)
   ,  CZI2  => c_z_int(1)
   ,  CZI3  => c_z_int(2)
   ,  CZI4  => c_z_int(3)
   ,  CZI5  => c_z_int(4)
   ,  CZI6  => c_z_int(5)
   ,  CZI7  => c_z_int(6)
   ,  CZI8  => c_z_int(7)
   ,  CZI9  => c_z_int(8)
   ,  CZI10 => c_z_int(9)
   ,  CZI11 => c_z_int(10)
   ,  CZI12 => c_z_int(11)
   ,  CZI13 => c_z_int(12)
   ,  CZI14 => c_z_int(13)
   ,  CZI15 => c_z_int(14)
   ,  CZI16 => c_z_int(15)
   ,  CZI17 => c_z_int(16)
   ,  CZI18 => c_z_int(17)
   ,  CZI19 => c_z_int(18)
   ,  CZI20 => c_z_int(19)
   ,  CZI21 => c_z_int(20)
   ,  CZI22 => c_z_int(21)
   ,  CZI23 => c_z_int(22)
   ,  CZI24 => c_z_int(23)
   ,  CZI25 => c_z_int(24)
   ,  CZI26 => c_z_int(25)
   ,  CZI27 => c_z_int(26)
   ,  CZI28 => c_z_int(27)
   ,  CZI29 => c_z_int(28)
   ,  CZI30 => c_z_int(29)
   ,  CZI31 => c_z_int(30)
   ,  CZI32 => c_z_int(31)
   ,  CZI33 => c_z_int(32)
   ,  CZI34 => c_z_int(33)
   ,  CZI35 => c_z_int(34)
   ,  CZI36 => c_z_int(35)
   ,  CZI37 => c_z_int(36)
   ,  CZI38 => c_z_int(37)
   ,  CZI39 => c_z_int(38)
   ,  CZI40 => c_z_int(39)
   ,  CZI41 => c_z_int(40)
   ,  CZI42 => c_z_int(41)
   ,  CZI43 => c_z_int(42)
   ,  CZI44 => c_z_int(43)
   ,  CZI45 => c_z_int(44)
   ,  CZI46 => c_z_int(45)
   ,  CZI47 => c_z_int(46)
   ,  CZI48 => c_z_int(47)
   ,  CZI49 => c_z_int(48)
   ,  CZI50 => c_z_int(49)
   ,  CZI51 => c_z_int(50)
   ,  CZI52 => c_z_int(51)
   ,  CZI53 => c_z_int(52)
   ,  CZI54 => c_z_int(53)
   ,  CZI55 => c_z_int(54)
   ,  CZI56 => c_z_int(55)
   ,  CZO1  => OPEN
   ,  CZO2  => OPEN
   ,  CZO3  => OPEN
   ,  CZO4  => OPEN
   ,  CZO5  => OPEN
   ,  CZO6  => OPEN
   ,  CZO7  => OPEN
   ,  CZO8  => OPEN
   ,  CZO9  => OPEN
   ,  CZO10 => OPEN
   ,  CZO11 => OPEN
   ,  CZO12 => OPEN
   ,  CZO13 => OPEN
   ,  CZO14 => OPEN
   ,  CZO15 => OPEN
   ,  CZO16 => OPEN
   ,  CZO17 => OPEN
   ,  CZO18 => OPEN
   ,  CZO19 => OPEN
   ,  CZO20 => OPEN
   ,  CZO21 => OPEN
   ,  CZO22 => OPEN
   ,  CZO23 => OPEN
   ,  CZO24 => OPEN
   ,  CZO25 => OPEN
   ,  CZO26 => OPEN
   ,  CZO27 => OPEN
   ,  CZO28 => OPEN
   ,  CZO29 => OPEN
   ,  CZO30 => OPEN
   ,  CZO31 => OPEN
   ,  CZO32 => OPEN
   ,  CZO33 => OPEN
   ,  CZO34 => OPEN
   ,  CZO35 => OPEN
   ,  CZO36 => OPEN
   ,  CZO37 => OPEN
   ,  CZO38 => OPEN
   ,  CZO39 => OPEN
   ,  CZO40 => OPEN
   ,  CZO41 => OPEN
   ,  CZO42 => OPEN
   ,  CZO43 => OPEN
   ,  CZO44 => OPEN
   ,  CZO45 => OPEN
   ,  CZO46 => OPEN
   ,  CZO47 => OPEN
   ,  CZO48 => OPEN
   ,  CZO49 => OPEN
   ,  CZO50 => OPEN
   ,  CZO51 => OPEN
   ,  CZO52 => OPEN
   ,  CZO53 => OPEN
   ,  CZO54 => OPEN
   ,  CZO55 => OPEN
   ,  CZO56 => OPEN
   ,  D1    => dsp0_d_i(0)
   ,  D2    => dsp0_d_i(1)
   ,  D3    => dsp0_d_i(2)
   ,  D4    => dsp0_d_i(3)
   ,  D5    => dsp0_d_i(4)
   ,  D6    => dsp0_d_i(5)
   ,  D7    => dsp0_d_i(6)
   ,  D8    => dsp0_d_i(7)
   ,  D9    => dsp0_d_i(8)
   ,  D10   => dsp0_d_i(9)
   ,  D11   => dsp0_d_i(10)
   ,  D12   => dsp0_d_i(11)
   ,  D13   => dsp0_d_i(12)
   ,  D14   => dsp0_d_i(13)
   ,  D15   => dsp0_d_i(14)
   ,  D16   => dsp0_d_i(15)
   ,  D17   => dsp0_d_i(16)
   ,  D18   => dsp0_d_i(17)
   ,  OVF   => dsp0_ovf_o
   ,  R     => dsp0_rst_i
   ,  RZ    => dsp0_rstz_i
   ,  WE    => dsp0_we_i
   ,  WEZ   => dsp0_wez_i
   ,  Z1    => dsp0_z_o(0)
   ,  Z2    => dsp0_z_o(1)
   ,  Z3    => dsp0_z_o(2)
   ,  Z4    => dsp0_z_o(3)
   ,  Z5    => dsp0_z_o(4)
   ,  Z6    => dsp0_z_o(5)
   ,  Z7    => dsp0_z_o(6)
   ,  Z8    => dsp0_z_o(7)
   ,  Z9    => dsp0_z_o(8)
   ,  Z10   => dsp0_z_o(9)
   ,  Z11   => dsp0_z_o(10)
   ,  Z12   => dsp0_z_o(11)
   ,  Z13   => dsp0_z_o(12)
   ,  Z14   => dsp0_z_o(13)
   ,  Z15   => dsp0_z_o(14)
   ,  Z16   => dsp0_z_o(15)
   ,  Z17   => dsp0_z_o(16)
   ,  Z18   => dsp0_z_o(17)
   ,  Z19   => dsp0_z_o(18)
   ,  Z20   => dsp0_z_o(19)
   ,  Z21   => dsp0_z_o(20)
   ,  Z22   => dsp0_z_o(21)
   ,  Z23   => dsp0_z_o(22)
   ,  Z24   => dsp0_z_o(23)
   ,  Z25   => dsp0_z_o(24)
   ,  Z26   => dsp0_z_o(25)
   ,  Z27   => dsp0_z_o(26)
   ,  Z28   => dsp0_z_o(27)
   ,  Z29   => dsp0_z_o(28)
   ,  Z30   => dsp0_z_o(29)
   ,  Z31   => dsp0_z_o(30)
   ,  Z32   => dsp0_z_o(31)
   ,  Z33   => dsp0_z_o(32)
   ,  Z34   => dsp0_z_o(33)
   ,  Z35   => dsp0_z_o(34)
   ,  Z36   => dsp0_z_o(35)
   ,  Z37   => dsp0_z_o(36)
   ,  Z38   => dsp0_z_o(37)
   ,  Z39   => dsp0_z_o(38)
   ,  Z40   => dsp0_z_o(39)
   ,  Z41   => dsp0_z_o(40)
   ,  Z42   => dsp0_z_o(41)
   ,  Z43   => dsp0_z_o(42)
   ,  Z44   => dsp0_z_o(43)
   ,  Z45   => dsp0_z_o(44)
   ,  Z46   => dsp0_z_o(45)
   ,  Z47   => dsp0_z_o(46)
   ,  Z48   => dsp0_z_o(47)
   ,  Z49   => dsp0_z_o(48)
   ,  Z50   => dsp0_z_o(49)
   ,  Z51   => dsp0_z_o(50)
   ,  Z52   => dsp0_z_o(51)
   ,  Z53   => dsp0_z_o(52)
   ,  Z54   => dsp0_z_o(53)
   ,  Z55   => dsp0_z_o(54)
   ,  Z56   => dsp0_z_o(55)
);
--#}}}#

-- instance dsp1#{{{#
dsp_1 : NX_DSP_U_BOX
generic map (
    col    => col
  , row    => row
  , cfg_bot_i => cfg_bot_i
  , cfg_top_i => cfg_top_i
)
port map (
      A1    => dsp1_a_i(0)
   ,  A2    => dsp1_a_i(1)
   ,  A3    => dsp1_a_i(2)
   ,  A4    => dsp1_a_i(3)
   ,  A5    => dsp1_a_i(4)
   ,  A6    => dsp1_a_i(5)
   ,  A7    => dsp1_a_i(6)
   ,  A8    => dsp1_a_i(7)
   ,  A9    => dsp1_a_i(8)
   ,  A10   => dsp1_a_i(9)
   ,  A11   => dsp1_a_i(10)
   ,  A12   => dsp1_a_i(11)
   ,  A13   => dsp1_a_i(12)
   ,  A14   => dsp1_a_i(13)
   ,  A15   => dsp1_a_i(14)
   ,  A16   => dsp1_a_i(15)
   ,  A17   => dsp1_a_i(16)
   ,  A18   => dsp1_a_i(17)
   ,  A19   => dsp1_a_i(18)
   ,  A20   => dsp1_a_i(19)
   ,  A21   => dsp1_a_i(20)
   ,  A22   => dsp1_a_i(21)
   ,  A23   => dsp1_a_i(22)
   ,  A24   => dsp1_a_i(23)
   ,  B1    => dsp1_b_i(0)
   ,  B2    => dsp1_b_i(1)
   ,  B3    => dsp1_b_i(2)
   ,  B4    => dsp1_b_i(3)
   ,  B5    => dsp1_b_i(4)
   ,  B6    => dsp1_b_i(5)
   ,  B7    => dsp1_b_i(6)
   ,  B8    => dsp1_b_i(7)
   ,  B9    => dsp1_b_i(8)
   ,  B10   => dsp1_b_i(9)
   ,  B11   => dsp1_b_i(10)
   ,  B12   => dsp1_b_i(11)
   ,  B13   => dsp1_b_i(12)
   ,  B14   => dsp1_b_i(13)
   ,  B15   => dsp1_b_i(14)
   ,  B16   => dsp1_b_i(15)
   ,  B17   => dsp1_b_i(16)
   ,  B18   => dsp1_b_i(17)
   ,  C1    => dsp1_c_i(0)
   ,  C2    => dsp1_c_i(1)
   ,  C3    => dsp1_c_i(2)
   ,  C4    => dsp1_c_i(3)
   ,  C5    => dsp1_c_i(4)
   ,  C6    => dsp1_c_i(5)
   ,  C7    => dsp1_c_i(6)
   ,  C8    => dsp1_c_i(7)
   ,  C9    => dsp1_c_i(8)
   ,  C10   => dsp1_c_i(9)
   ,  C11   => dsp1_c_i(10)
   ,  C12   => dsp1_c_i(11)
   ,  C13   => dsp1_c_i(12)
   ,  C14   => dsp1_c_i(13)
   ,  C15   => dsp1_c_i(14)
   ,  C16   => dsp1_c_i(15)
   ,  C17   => dsp1_c_i(16)
   ,  C18   => dsp1_c_i(17)
   ,  C19   => dsp1_c_i(18)
   ,  C20   => dsp1_c_i(19)
   ,  C21   => dsp1_c_i(20)
   ,  C22   => dsp1_c_i(21)
   ,  C23   => dsp1_c_i(22)
   ,  C24   => dsp1_c_i(23)
   ,  C25   => dsp1_c_i(24)
   ,  C26   => dsp1_c_i(25)
   ,  C27   => dsp1_c_i(26)
   ,  C28   => dsp1_c_i(27)
   ,  C29   => dsp1_c_i(28)
   ,  C30   => dsp1_c_i(29)
   ,  C31   => dsp1_c_i(30)
   ,  C32   => dsp1_c_i(31)
   ,  C33   => dsp1_c_i(32)
   ,  C34   => dsp1_c_i(33)
   ,  C35   => dsp1_c_i(34)
   ,  C36   => dsp1_c_i(35)
   ,  CAI1  => '0'
   ,  CAI2  => '0'
   ,  CAI3  => '0'
   ,  CAI4  => '0'
   ,  CAI5  => '0'
   ,  CAI6  => '0'
   ,  CAI7  => '0'
   ,  CAI8  => '0'
   ,  CAI9  => '0'
   ,  CAI10 => '0'
   ,  CAI11 => '0'
   ,  CAI12 => '0'
   ,  CAI13 => '0'
   ,  CAI14 => '0'
   ,  CAI15 => '0'
   ,  CAI16 => '0'
   ,  CAI17 => '0'
   ,  CAI18 => '0'
   ,  CAI19 => '0'
   ,  CAI20 => '0'
   ,  CAI21 => '0'
   ,  CAI22 => '0'
   ,  CAI23 => '0'
   ,  CAI24 => '0'
   ,  CAO1  => c_a_int(0)
   ,  CAO2  => c_a_int(1)
   ,  CAO3  => c_a_int(2)
   ,  CAO4  => c_a_int(3)
   ,  CAO5  => c_a_int(4)
   ,  CAO6  => c_a_int(5)
   ,  CAO7  => c_a_int(6)
   ,  CAO8  => c_a_int(7)
   ,  CAO9  => c_a_int(8)
   ,  CAO10 => c_a_int(9)
   ,  CAO11 => c_a_int(10)
   ,  CAO12 => c_a_int(11)
   ,  CAO13 => c_a_int(12)
   ,  CAO14 => c_a_int(13)
   ,  CAO15 => c_a_int(14)
   ,  CAO16 => c_a_int(15)
   ,  CAO17 => c_a_int(16)
   ,  CAO18 => c_a_int(17)
   ,  CAO19 => c_a_int(18)
   ,  CAO20 => c_a_int(19)
   ,  CAO21 => c_a_int(20)
   ,  CAO22 => c_a_int(21)
   ,  CAO23 => c_a_int(22)
   ,  CAO24 => c_a_int(23)
   ,  CBI1  => '0'
   ,  CBI2  => '0'
   ,  CBI3  => '0'
   ,  CBI4  => '0'
   ,  CBI5  => '0'
   ,  CBI6  => '0'
   ,  CBI7  => '0'
   ,  CBI8  => '0'
   ,  CBI9  => '0'
   ,  CBI10 => '0'
   ,  CBI11 => '0'
   ,  CBI12 => '0'
   ,  CBI13 => '0'
   ,  CBI14 => '0'
   ,  CBI15 => '0'
   ,  CBI16 => '0'
   ,  CBI17 => '0'
   ,  CBI18 => '0'
   ,  CBO1  => c_b_int(0)
   ,  CBO2  => c_b_int(1)
   ,  CBO3  => c_b_int(2)
   ,  CBO4  => c_b_int(3)
   ,  CBO5  => c_b_int(4)
   ,  CBO6  => c_b_int(5)
   ,  CBO7  => c_b_int(6)
   ,  CBO8  => c_b_int(7)
   ,  CBO9  => c_b_int(8)
   ,  CBO10 => c_b_int(9)
   ,  CBO11 => c_b_int(10)
   ,  CBO12 => c_b_int(11)
   ,  CBO13 => c_b_int(12)
   ,  CBO14 => c_b_int(13)
   ,  CBO15 => c_b_int(14)
   ,  CBO16 => c_b_int(15)
   ,  CBO17 => c_b_int(16)
   ,  CBO18 => c_b_int(17)
   ,  CCI   => c_cy_int
   ,  CCO   => OPEN
   ,  CI    => dsp1_cy_i
   ,  CK    => dsp1_clk_i
   ,  RESERVED => dsp1_cy_o
   ,  CO43  => dsp1_cy42_o
   ,  CO57  => dsp1_cy56_o
   ,  CZI1  => '0'
   ,  CZI2  => '0'
   ,  CZI3  => '0'
   ,  CZI4  => '0'
   ,  CZI5  => '0'
   ,  CZI6  => '0'
   ,  CZI7  => '0'
   ,  CZI8  => '0'
   ,  CZI9  => '0'
   ,  CZI10 => '0'
   ,  CZI11 => '0'
   ,  CZI12 => '0'
   ,  CZI13 => '0'
   ,  CZI14 => '0'
   ,  CZI15 => '0'
   ,  CZI16 => '0'
   ,  CZI17 => '0'
   ,  CZI18 => '0'
   ,  CZI19 => '0'
   ,  CZI20 => '0'
   ,  CZI21 => '0'
   ,  CZI22 => '0'
   ,  CZI23 => '0'
   ,  CZI24 => '0'
   ,  CZI25 => '0'
   ,  CZI26 => '0'
   ,  CZI27 => '0'
   ,  CZI28 => '0'
   ,  CZI29 => '0'
   ,  CZI30 => '0'
   ,  CZI31 => '0'
   ,  CZI32 => '0'
   ,  CZI33 => '0'
   ,  CZI34 => '0'
   ,  CZI35 => '0'
   ,  CZI36 => '0'
   ,  CZI37 => '0'
   ,  CZI38 => '0'
   ,  CZI39 => '0'
   ,  CZI40 => '0'
   ,  CZI41 => '0'
   ,  CZI42 => '0'
   ,  CZI43 => '0'
   ,  CZI44 => '0'
   ,  CZI45 => '0'
   ,  CZI46 => '0'
   ,  CZI47 => '0'
   ,  CZI48 => '0'
   ,  CZI49 => '0'
   ,  CZI50 => '0'
   ,  CZI51 => '0'
   ,  CZI52 => '0'
   ,  CZI53 => '0'
   ,  CZI54 => '0'
   ,  CZI55 => '0'
   ,  CZI56 => '0'
   ,  CZO1  => c_z_int(0)
   ,  CZO2  => c_z_int(1)
   ,  CZO3  => c_z_int(2)
   ,  CZO4  => c_z_int(3)
   ,  CZO5  => c_z_int(4)
   ,  CZO6  => c_z_int(5)
   ,  CZO7  => c_z_int(6)
   ,  CZO8  => c_z_int(7)
   ,  CZO9  => c_z_int(8)
   ,  CZO10 => c_z_int(9)
   ,  CZO11 => c_z_int(10)
   ,  CZO12 => c_z_int(11)
   ,  CZO13 => c_z_int(12)
   ,  CZO14 => c_z_int(13)
   ,  CZO15 => c_z_int(14)
   ,  CZO16 => c_z_int(15)
   ,  CZO17 => c_z_int(16)
   ,  CZO18 => c_z_int(17)
   ,  CZO19 => c_z_int(18)
   ,  CZO20 => c_z_int(19)
   ,  CZO21 => c_z_int(20)
   ,  CZO22 => c_z_int(21)
   ,  CZO23 => c_z_int(22)
   ,  CZO24 => c_z_int(23)
   ,  CZO25 => c_z_int(24)
   ,  CZO26 => c_z_int(25)
   ,  CZO27 => c_z_int(26)
   ,  CZO28 => c_z_int(27)
   ,  CZO29 => c_z_int(28)
   ,  CZO30 => c_z_int(29)
   ,  CZO31 => c_z_int(30)
   ,  CZO32 => c_z_int(31)
   ,  CZO33 => c_z_int(32)
   ,  CZO34 => c_z_int(33)
   ,  CZO35 => c_z_int(34)
   ,  CZO36 => c_z_int(35)
   ,  CZO37 => c_z_int(36)
   ,  CZO38 => c_z_int(37)
   ,  CZO39 => c_z_int(38)
   ,  CZO40 => c_z_int(39)
   ,  CZO41 => c_z_int(40)
   ,  CZO42 => c_z_int(41)
   ,  CZO43 => c_z_int(42)
   ,  CZO44 => c_z_int(43)
   ,  CZO45 => c_z_int(44)
   ,  CZO46 => c_z_int(45)
   ,  CZO47 => c_z_int(46)
   ,  CZO48 => c_z_int(47)
   ,  CZO49 => c_z_int(48)
   ,  CZO50 => c_z_int(49)
   ,  CZO51 => c_z_int(50)
   ,  CZO52 => c_z_int(51)
   ,  CZO53 => c_z_int(52)
   ,  CZO54 => c_z_int(53)
   ,  CZO55 => c_z_int(54)
   ,  CZO56 => c_z_int(55)
   ,  D1    => dsp1_d_i(0)
   ,  D2    => dsp1_d_i(1)
   ,  D3    => dsp1_d_i(2)
   ,  D4    => dsp1_d_i(3)
   ,  D5    => dsp1_d_i(4)
   ,  D6    => dsp1_d_i(5)
   ,  D7    => dsp1_d_i(6)
   ,  D8    => dsp1_d_i(7)
   ,  D9    => dsp1_d_i(8)
   ,  D10   => dsp1_d_i(9)
   ,  D11   => dsp1_d_i(10)
   ,  D12   => dsp1_d_i(11)
   ,  D13   => dsp1_d_i(12)
   ,  D14   => dsp1_d_i(13)
   ,  D15   => dsp1_d_i(14)
   ,  D16   => dsp1_d_i(15)
   ,  D17   => dsp1_d_i(16)
   ,  D18   => dsp1_d_i(17)
   ,  OVF   => dsp1_ovf_o
   ,  R     => dsp1_rst_i
   ,  RZ    => dsp1_rstz_i
   ,  WE    => dsp1_we_i
   ,  WEZ   => dsp1_wez_i
   ,  Z1    => dsp1_z_o(0)
   ,  Z2    => dsp1_z_o(1)
   ,  Z3    => dsp1_z_o(2)
   ,  Z4    => dsp1_z_o(3)
   ,  Z5    => dsp1_z_o(4)
   ,  Z6    => dsp1_z_o(5)
   ,  Z7    => dsp1_z_o(6)
   ,  Z8    => dsp1_z_o(7)
   ,  Z9    => dsp1_z_o(8)
   ,  Z10   => dsp1_z_o(9)
   ,  Z11   => dsp1_z_o(10)
   ,  Z12   => dsp1_z_o(11)
   ,  Z13   => dsp1_z_o(12)
   ,  Z14   => dsp1_z_o(13)
   ,  Z15   => dsp1_z_o(14)
   ,  Z16   => dsp1_z_o(15)
   ,  Z17   => dsp1_z_o(16)
   ,  Z18   => dsp1_z_o(17)
   ,  Z19   => dsp1_z_o(18)
   ,  Z20   => dsp1_z_o(19)
   ,  Z21   => dsp1_z_o(20)
   ,  Z22   => dsp1_z_o(21)
   ,  Z23   => dsp1_z_o(22)
   ,  Z24   => dsp1_z_o(23)
   ,  Z25   => dsp1_z_o(24)
   ,  Z26   => dsp1_z_o(25)
   ,  Z27   => dsp1_z_o(26)
   ,  Z28   => dsp1_z_o(27)
   ,  Z29   => dsp1_z_o(28)
   ,  Z30   => dsp1_z_o(29)
   ,  Z31   => dsp1_z_o(30)
   ,  Z32   => dsp1_z_o(31)
   ,  Z33   => dsp1_z_o(32)
   ,  Z34   => dsp1_z_o(33)
   ,  Z35   => dsp1_z_o(34)
   ,  Z36   => dsp1_z_o(35)
   ,  Z37   => dsp1_z_o(36)
   ,  Z38   => dsp1_z_o(37)
   ,  Z39   => dsp1_z_o(38)
   ,  Z40   => dsp1_z_o(39)
   ,  Z41   => dsp1_z_o(40)
   ,  Z42   => dsp1_z_o(41)
   ,  Z43   => dsp1_z_o(42)
   ,  Z44   => dsp1_z_o(43)
   ,  Z45   => dsp1_z_o(44)
   ,  Z46   => dsp1_z_o(45)
   ,  Z47   => dsp1_z_o(46)
   ,  Z48   => dsp1_z_o(47)
   ,  Z49   => dsp1_z_o(48)
   ,  Z50   => dsp1_z_o(49)
   ,  Z51   => dsp1_z_o(50)
   ,  Z52   => dsp1_z_o(51)
   ,  Z53   => dsp1_z_o(52)
   ,  Z54   => dsp1_z_o(53)
   ,  Z55   => dsp1_z_o(54)
   ,  Z56   => dsp1_z_o(55)
);
--#}}}#

-- instance ram0#{{{#
ram_0 : NX_RAM_U_BOX
generic map (
    col    => col
  , row    => row
  , cfg_bot_i => cfg_bot_i
  , cfg_top_i => cfg_top_i
)
port map (
    ACK   => dpram_clkmem0_i
  , BCK   => dpram_clkmem1_i

  , AI1   => dpram_din0_i(0)
  , AI2   => dpram_din0_i(1)
  , AI3   => dpram_din0_i(2)
  , AI4   => dpram_din0_i(3)
  , AI5   => dpram_din0_i(4)
  , AI6   => dpram_din0_i(5)
  , AI7   => dpram_din0_i(6)
  , AI8   => dpram_din0_i(7)
  , AI9   => dpram_din0_i(8)
  , AI10  => dpram_din0_i(9)
  , AI11  => dpram_din0_i(10)
  , AI12  => dpram_din0_i(11)
  , AI13  => dpram_din0_i(12)
  , AI14  => dpram_din0_i(13)
  , AI15  => dpram_din0_i(14)
  , AI16  => dpram_din0_i(15)
  , AI17  => dpram_din0_i(16)
  , AI18  => dpram_din0_i(17)
  , AI19  => dpram_din0_i(18)
  , AI20  => dpram_din0_i(19)
  , AI21  => dpram_din0_i(20)
  , AI22  => dpram_din0_i(21)
  , AI23  => dpram_din0_i(22)
  , AI24  => dpram_din0_i(23)

  , BI1   => dpram_din1_i(0)
  , BI2   => dpram_din1_i(1)
  , BI3   => dpram_din1_i(2)
  , BI4   => dpram_din1_i(3)
  , BI5   => dpram_din1_i(4)
  , BI6   => dpram_din1_i(5)
  , BI7   => dpram_din1_i(6)
  , BI8   => dpram_din1_i(7)
  , BI9   => dpram_din1_i(8)
  , BI10  => dpram_din1_i(9)
  , BI11  => dpram_din1_i(10)
  , BI12  => dpram_din1_i(11)
  , BI13  => dpram_din1_i(12)
  , BI14  => dpram_din1_i(13)
  , BI15  => dpram_din1_i(14)
  , BI16  => dpram_din1_i(15)
  , BI17  => dpram_din1_i(16)
  , BI18  => dpram_din1_i(17)
  , BI19  => dpram_din1_i(18)
  , BI20  => dpram_din1_i(19)
  , BI21  => dpram_din1_i(20)
  , BI22  => dpram_din1_i(21)
  , BI23  => dpram_din1_i(22)
  , BI24  => dpram_din1_i(23)

  , ACOR => dpram_ecc_corrected0_o
  , AERR => dpram_ecc_uncorrected0_o
  , BCOR => dpram_ecc_corrected1_o
  , BERR => dpram_ecc_uncorrected1_o

  , AO1  => dpram_dout0_o(0)
  , AO2  => dpram_dout0_o(1)
  , AO3  => dpram_dout0_o(2)
  , AO4  => dpram_dout0_o(3)
  , AO5  => dpram_dout0_o(4)
  , AO6  => dpram_dout0_o(5)
  , AO7  => dpram_dout0_o(6)
  , AO8  => dpram_dout0_o(7)
  , AO9  => dpram_dout0_o(8)
  , AO10 => dpram_dout0_o(9)
  , AO11 => dpram_dout0_o(10)
  , AO12 => dpram_dout0_o(11)
  , AO13 => dpram_dout0_o(12)
  , AO14 => dpram_dout0_o(13)
  , AO15 => dpram_dout0_o(14)
  , AO16 => dpram_dout0_o(15)
  , AO17 => dpram_dout0_o(16)
  , AO18 => dpram_dout0_o(17)
  , AO19 => dpram_dout0_o(18)
  , AO20 => dpram_dout0_o(19)
  , AO21 => dpram_dout0_o(20)
  , AO22 => dpram_dout0_o(21)
  , AO23 => dpram_dout0_o(22)
  , AO24 => dpram_dout0_o(23)

  , BO1  => dpram_dout1_o(0)
  , BO2  => dpram_dout1_o(1)
  , BO3  => dpram_dout1_o(2)
  , BO4  => dpram_dout1_o(3)
  , BO5  => dpram_dout1_o(4)
  , BO6  => dpram_dout1_o(5)
  , BO7  => dpram_dout1_o(6)
  , BO8  => dpram_dout1_o(7)
  , BO9  => dpram_dout1_o(8)
  , BO10 => dpram_dout1_o(9)
  , BO11 => dpram_dout1_o(10)
  , BO12 => dpram_dout1_o(11)
  , BO13 => dpram_dout1_o(12)
  , BO14 => dpram_dout1_o(13)
  , BO15 => dpram_dout1_o(14)
  , BO16 => dpram_dout1_o(15)
  , BO17 => dpram_dout1_o(16)
  , BO18 => dpram_dout1_o(17)
  , BO19 => dpram_dout1_o(18)
  , BO20 => dpram_dout1_o(19)
  , BO21 => dpram_dout1_o(20)
  , BO22 => dpram_dout1_o(21)
  , BO23 => dpram_dout1_o(22)
  , BO24 => dpram_dout1_o(23)

  , AA1  => dpram_addr0_i(0)
  , AA2  => dpram_addr0_i(1)
  , AA3  => dpram_addr0_i(2)
  , AA4  => dpram_addr0_i(3)
  , AA5  => dpram_addr0_i(4)
  , AA6  => dpram_addr0_i(5)
  , AA7  => dpram_addr0_i(6)
  , AA8  => dpram_addr0_i(7)
  , AA9  => dpram_addr0_i(8)
  , AA10 => dpram_addr0_i(9)
  , AA11 => dpram_addr0_i(10)
  , AA12 => dpram_addr0_i(11)
  , AA13 => dpram_addr0_i(12)
  , AA14 => dpram_addr0_i(13)
  , AA15 => dpram_addr0_i(14)
  , AA16 => dpram_addr0_i(15)

  , ACS  => dpram_cs0_i
  , AWE  => dpram_we0_i
  , AR   => dpram_rst0_i

  , BA1  => dpram_addr1_i(0)
  , BA2  => dpram_addr1_i(1)
  , BA3  => dpram_addr1_i(2)
  , BA4  => dpram_addr1_i(3)
  , BA5  => dpram_addr1_i(4)
  , BA6  => dpram_addr1_i(5)
  , BA7  => dpram_addr1_i(6)
  , BA8  => dpram_addr1_i(7)
  , BA9  => dpram_addr1_i(8)
  , BA10 => dpram_addr1_i(9)
  , BA11 => dpram_addr1_i(10)
  , BA12 => dpram_addr1_i(11)
  , BA13 => dpram_addr1_i(12)
  , BA14 => dpram_addr1_i(13)
  , BA15 => dpram_addr1_i(14)
  , BA16 => dpram_addr1_i(15)

  , BCS  => dpram_cs1_i
  , BWE  => dpram_we1_i
  , BR   => dpram_rst1_i
);
--#}}}#

end NX_RTL;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_U_BOX definition
-- =================================================================================================

-- NX_DSP_U_BOX#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_DSP_U_BOX is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    A1    : in  std_logic;
    A2    : in  std_logic;
    A3    : in  std_logic;
    A4    : in  std_logic;
    A5    : in  std_logic;
    A6    : in  std_logic;
    A7    : in  std_logic;
    A8    : in  std_logic;
    A9    : in  std_logic;
    A10   : in  std_logic;
    A11   : in  std_logic;
    A12   : in  std_logic;
    A13   : in  std_logic;
    A14   : in  std_logic;
    A15   : in  std_logic;
    A16   : in  std_logic;
    A17   : in  std_logic;
    A18   : in  std_logic;
    A19   : in  std_logic;
    A20   : in  std_logic;
    A21   : in  std_logic;
    A22   : in  std_logic;
    A23   : in  std_logic;
    A24   : in  std_logic;

    B1    : in  std_logic;
    B2    : in  std_logic;
    B3    : in  std_logic;
    B4    : in  std_logic;
    B5    : in  std_logic;
    B6    : in  std_logic;
    B7    : in  std_logic;
    B8    : in  std_logic;
    B9    : in  std_logic;
    B10   : in  std_logic;
    B11   : in  std_logic;
    B12   : in  std_logic;
    B13   : in  std_logic;
    B14   : in  std_logic;
    B15   : in  std_logic;
    B16   : in  std_logic;
    B17   : in  std_logic;
    B18   : in  std_logic;

    C1    : in  std_logic;
    C2    : in  std_logic;
    C3    : in  std_logic;
    C4    : in  std_logic;
    C5    : in  std_logic;
    C6    : in  std_logic;
    C7    : in  std_logic;
    C8    : in  std_logic;
    C9    : in  std_logic;
    C10   : in  std_logic;
    C11   : in  std_logic;
    C12   : in  std_logic;
    C13   : in  std_logic;
    C14   : in  std_logic;
    C15   : in  std_logic;
    C16   : in  std_logic;
    C17   : in  std_logic;
    C18   : in  std_logic;
    C19   : in  std_logic;
    C20   : in  std_logic;
    C21   : in  std_logic;
    C22   : in  std_logic;
    C23   : in  std_logic;
    C24   : in  std_logic;
    C25   : in  std_logic;
    C26   : in  std_logic;
    C27   : in  std_logic;
    C28   : in  std_logic;
    C29   : in  std_logic;
    C30   : in  std_logic;
    C31   : in  std_logic;
    C32   : in  std_logic;
    C33   : in  std_logic;
    C34   : in  std_logic;
    C35   : in  std_logic;
    C36   : in  std_logic;

    CAI1  : in  std_logic;
    CAI2  : in  std_logic;
    CAI3  : in  std_logic;
    CAI4  : in  std_logic;
    CAI5  : in  std_logic;
    CAI6  : in  std_logic;
    CAI7  : in  std_logic;
    CAI8  : in  std_logic;
    CAI9  : in  std_logic;
    CAI10 : in  std_logic;
    CAI11 : in  std_logic;
    CAI12 : in  std_logic;
    CAI13 : in  std_logic;
    CAI14 : in  std_logic;
    CAI15 : in  std_logic;
    CAI16 : in  std_logic;
    CAI17 : in  std_logic;
    CAI18 : in  std_logic;
    CAI19 : in  std_logic;
    CAI20 : in  std_logic;
    CAI21 : in  std_logic;
    CAI22 : in  std_logic;
    CAI23 : in  std_logic;
    CAI24 : in  std_logic;

    CAO1  : out std_logic;
    CAO2  : out std_logic;
    CAO3  : out std_logic;
    CAO4  : out std_logic;
    CAO5  : out std_logic;
    CAO6  : out std_logic;
    CAO7  : out std_logic;
    CAO8  : out std_logic;
    CAO9  : out std_logic;
    CAO10 : out std_logic;
    CAO11 : out std_logic;
    CAO12 : out std_logic;
    CAO13 : out std_logic;
    CAO14 : out std_logic;
    CAO15 : out std_logic;
    CAO16 : out std_logic;
    CAO17 : out std_logic;
    CAO18 : out std_logic;
    CAO19 : out std_logic;
    CAO20 : out std_logic;
    CAO21 : out std_logic;
    CAO22 : out std_logic;
    CAO23 : out std_logic;
    CAO24 : out std_logic;

    CBI1  : in  std_logic;
    CBI2  : in  std_logic;
    CBI3  : in  std_logic;
    CBI4  : in  std_logic;
    CBI5  : in  std_logic;
    CBI6  : in  std_logic;
    CBI7  : in  std_logic;
    CBI8  : in  std_logic;
    CBI9  : in  std_logic;
    CBI10 : in  std_logic;
    CBI11 : in  std_logic;
    CBI12 : in  std_logic;
    CBI13 : in  std_logic;
    CBI14 : in  std_logic;
    CBI15 : in  std_logic;
    CBI16 : in  std_logic;
    CBI17 : in  std_logic;
    CBI18 : in  std_logic;

    CBO1  : out std_logic;
    CBO2  : out std_logic;
    CBO3  : out std_logic;
    CBO4  : out std_logic;
    CBO5  : out std_logic;
    CBO6  : out std_logic;
    CBO7  : out std_logic;
    CBO8  : out std_logic;
    CBO9  : out std_logic;
    CBO10 : out std_logic;
    CBO11 : out std_logic;
    CBO12 : out std_logic;
    CBO13 : out std_logic;
    CBO14 : out std_logic;
    CBO15 : out std_logic;
    CBO16 : out std_logic;
    CBO17 : out std_logic;
    CBO18 : out std_logic;

    CCI   : in  std_logic;
    CCO   : out std_logic;
    CI    : in  std_logic;
    CK    : in  std_logic;
    RESERVED: out std_logic;
    CO43  : out std_logic;
    CO57  : out std_logic;

    CZI1  : in  std_logic;
    CZI2  : in  std_logic;
    CZI3  : in  std_logic;
    CZI4  : in  std_logic;
    CZI5  : in  std_logic;
    CZI6  : in  std_logic;
    CZI7  : in  std_logic;
    CZI8  : in  std_logic;
    CZI9  : in  std_logic;
    CZI10 : in  std_logic;
    CZI11 : in  std_logic;
    CZI12 : in  std_logic;
    CZI13 : in  std_logic;
    CZI14 : in  std_logic;
    CZI15 : in  std_logic;
    CZI16 : in  std_logic;
    CZI17 : in  std_logic;
    CZI18 : in  std_logic;
    CZI19 : in  std_logic;
    CZI20 : in  std_logic;
    CZI21 : in  std_logic;
    CZI22 : in  std_logic;
    CZI23 : in  std_logic;
    CZI24 : in  std_logic;
    CZI25 : in  std_logic;
    CZI26 : in  std_logic;
    CZI27 : in  std_logic;
    CZI28 : in  std_logic;
    CZI29 : in  std_logic;
    CZI30 : in  std_logic;
    CZI31 : in  std_logic;
    CZI32 : in  std_logic;
    CZI33 : in  std_logic;
    CZI34 : in  std_logic;
    CZI35 : in  std_logic;
    CZI36 : in  std_logic;
    CZI37 : in  std_logic;
    CZI38 : in  std_logic;
    CZI39 : in  std_logic;
    CZI40 : in  std_logic;
    CZI41 : in  std_logic;
    CZI42 : in  std_logic;
    CZI43 : in  std_logic;
    CZI44 : in  std_logic;
    CZI45 : in  std_logic;
    CZI46 : in  std_logic;
    CZI47 : in  std_logic;
    CZI48 : in  std_logic;
    CZI49 : in  std_logic;
    CZI50 : in  std_logic;
    CZI51 : in  std_logic;
    CZI52 : in  std_logic;
    CZI53 : in  std_logic;
    CZI54 : in  std_logic;
    CZI55 : in  std_logic;
    CZI56 : in  std_logic;

    CZO1  : out std_logic;
    CZO2  : out std_logic;
    CZO3  : out std_logic;
    CZO4  : out std_logic;
    CZO5  : out std_logic;
    CZO6  : out std_logic;
    CZO7  : out std_logic;
    CZO8  : out std_logic;
    CZO9  : out std_logic;
    CZO10 : out std_logic;
    CZO11 : out std_logic;
    CZO12 : out std_logic;
    CZO13 : out std_logic;
    CZO14 : out std_logic;
    CZO15 : out std_logic;
    CZO16 : out std_logic;
    CZO17 : out std_logic;
    CZO18 : out std_logic;
    CZO19 : out std_logic;
    CZO20 : out std_logic;
    CZO21 : out std_logic;
    CZO22 : out std_logic;
    CZO23 : out std_logic;
    CZO24 : out std_logic;
    CZO25 : out std_logic;
    CZO26 : out std_logic;
    CZO27 : out std_logic;
    CZO28 : out std_logic;
    CZO29 : out std_logic;
    CZO30 : out std_logic;
    CZO31 : out std_logic;
    CZO32 : out std_logic;
    CZO33 : out std_logic;
    CZO34 : out std_logic;
    CZO35 : out std_logic;
    CZO36 : out std_logic;
    CZO37 : out std_logic;
    CZO38 : out std_logic;
    CZO39 : out std_logic;
    CZO40 : out std_logic;
    CZO41 : out std_logic;
    CZO42 : out std_logic;
    CZO43 : out std_logic;
    CZO44 : out std_logic;
    CZO45 : out std_logic;
    CZO46 : out std_logic;
    CZO47 : out std_logic;
    CZO48 : out std_logic;
    CZO49 : out std_logic;
    CZO50 : out std_logic;
    CZO51 : out std_logic;
    CZO52 : out std_logic;
    CZO53 : out std_logic;
    CZO54 : out std_logic;
    CZO55 : out std_logic;
    CZO56 : out std_logic;

    D1    : in  std_logic;
    D2    : in  std_logic;
    D3    : in  std_logic;
    D4    : in  std_logic;
    D5    : in  std_logic;
    D6    : in  std_logic;
    D7    : in  std_logic;
    D8    : in  std_logic;
    D9    : in  std_logic;
    D10   : in  std_logic;
    D11   : in  std_logic;
    D12   : in  std_logic;
    D13   : in  std_logic;
    D14   : in  std_logic;
    D15   : in  std_logic;
    D16   : in  std_logic;
    D17   : in  std_logic;
    D18   : in  std_logic;

    OVF   : out std_logic;
    R     : in  std_logic;
    RZ    : in  std_logic;
    WE    : in  std_logic;
    WEZ   : in  std_logic;

    Z1    : out std_logic;
    Z2    : out std_logic;
    Z3    : out std_logic;
    Z4    : out std_logic;
    Z5    : out std_logic;
    Z6    : out std_logic;
    Z7    : out std_logic;
    Z8    : out std_logic;
    Z9    : out std_logic;
    Z10   : out std_logic;
    Z11   : out std_logic;
    Z12   : out std_logic;
    Z13   : out std_logic;
    Z14   : out std_logic;
    Z15   : out std_logic;
    Z16   : out std_logic;
    Z17   : out std_logic;
    Z18   : out std_logic;
    Z19   : out std_logic;
    Z20   : out std_logic;
    Z21   : out std_logic;
    Z22   : out std_logic;
    Z23   : out std_logic;
    Z24   : out std_logic;
    Z25   : out std_logic;
    Z26   : out std_logic;
    Z27   : out std_logic;
    Z28   : out std_logic;
    Z29   : out std_logic;
    Z30   : out std_logic;
    Z31   : out std_logic;
    Z32   : out std_logic;
    Z33   : out std_logic;
    Z34   : out std_logic;
    Z35   : out std_logic;
    Z36   : out std_logic;
    Z37   : out std_logic;
    Z38   : out std_logic;
    Z39   : out std_logic;
    Z40   : out std_logic;
    Z41   : out std_logic;
    Z42   : out std_logic;
    Z43   : out std_logic;
    Z44   : out std_logic;
    Z45   : out std_logic;
    Z46   : out std_logic;
    Z47   : out std_logic;
    Z48   : out std_logic;
    Z49   : out std_logic;
    Z50   : out std_logic;
    Z51   : out std_logic;
    Z52   : out std_logic;
    Z53   : out std_logic;
    Z54   : out std_logic;
    Z55   : out std_logic;
    Z56   : out std_logic
);
end NX_DSP_U_BOX;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RAM_U_BOX definition
-- =================================================================================================

-- NX_RAM_U_BOX #{{{#
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_RAM_U_BOX is
generic (
    col    : integer := 2;
    row    : integer := 6;
    cfg_bot_i : bit_vector(95 downto 0) := (others => '0');
    cfg_top_i : bit_vector(95 downto 0) := (others => '0')
);
port (
    ACK   : in  std_logic;
    BCK   : in  std_logic;

    AI1   : in  std_logic;
    AI2   : in  std_logic;
    AI3   : in  std_logic;
    AI4   : in  std_logic;
    AI5   : in  std_logic;
    AI6   : in  std_logic;
    AI7   : in  std_logic;
    AI8   : in  std_logic;
    AI9   : in  std_logic;
    AI10  : in  std_logic;
    AI11  : in  std_logic;
    AI12  : in  std_logic;
    AI13  : in  std_logic;
    AI14  : in  std_logic;
    AI15  : in  std_logic;
    AI16  : in  std_logic;
    AI17  : in  std_logic;
    AI18  : in  std_logic;
    AI19  : in  std_logic;
    AI20  : in  std_logic;
    AI21  : in  std_logic;
    AI22  : in  std_logic;
    AI23  : in  std_logic;
    AI24  : in  std_logic;

    BI1   : in  std_logic;
    BI2   : in  std_logic;
    BI3   : in  std_logic;
    BI4   : in  std_logic;
    BI5   : in  std_logic;
    BI6   : in  std_logic;
    BI7   : in  std_logic;
    BI8   : in  std_logic;
    BI9   : in  std_logic;
    BI10  : in  std_logic;
    BI11  : in  std_logic;
    BI12  : in  std_logic;
    BI13  : in  std_logic;
    BI14  : in  std_logic;
    BI15  : in  std_logic;
    BI16  : in  std_logic;
    BI17  : in  std_logic;
    BI18  : in  std_logic;
    BI19  : in  std_logic;
    BI20  : in  std_logic;
    BI21  : in  std_logic;
    BI22  : in  std_logic;
    BI23  : in  std_logic;
    BI24  : in  std_logic;

    ACOR  : out std_logic;
    AERR  : out std_logic;
    BCOR  : out std_logic;
    BERR  : out std_logic;

    AO1   : out std_logic;
    AO2   : out std_logic;
    AO3   : out std_logic;
    AO4   : out std_logic;
    AO5   : out std_logic;
    AO6   : out std_logic;
    AO7   : out std_logic;
    AO8   : out std_logic;
    AO9   : out std_logic;
    AO10  : out std_logic;
    AO11  : out std_logic;
    AO12  : out std_logic;
    AO13  : out std_logic;
    AO14  : out std_logic;
    AO15  : out std_logic;
    AO16  : out std_logic;
    AO17  : out std_logic;
    AO18  : out std_logic;
    AO19  : out std_logic;
    AO20  : out std_logic;
    AO21  : out std_logic;
    AO22  : out std_logic;
    AO23  : out std_logic;
    AO24  : out std_logic;

    BO1   : out std_logic;
    BO2   : out std_logic;
    BO3   : out std_logic;
    BO4   : out std_logic;
    BO5   : out std_logic;
    BO6   : out std_logic;
    BO7   : out std_logic;
    BO8   : out std_logic;
    BO9   : out std_logic;
    BO10  : out std_logic;
    BO11  : out std_logic;
    BO12  : out std_logic;
    BO13  : out std_logic;
    BO14  : out std_logic;
    BO15  : out std_logic;
    BO16  : out std_logic;
    BO17  : out std_logic;
    BO18  : out std_logic;
    BO19  : out std_logic;
    BO20  : out std_logic;
    BO21  : out std_logic;
    BO22  : out std_logic;
    BO23  : out std_logic;
    BO24  : out std_logic;

    AA1   : in  std_logic;
    AA2   : in  std_logic;
    AA3   : in  std_logic;
    AA4   : in  std_logic;
    AA5   : in  std_logic;
    AA6   : in  std_logic;
    AA7   : in  std_logic;
    AA8   : in  std_logic;
    AA9   : in  std_logic;
    AA10  : in  std_logic;
    AA11  : in  std_logic;
    AA12  : in  std_logic;
    AA13  : in  std_logic;
    AA14  : in  std_logic;
    AA15  : in  std_logic;
    AA16  : in  std_logic;

    ACS   : in  std_logic;
    AWE   : in  std_logic;
    AR    : in  std_logic;

    BA1   : in  std_logic;
    BA2   : in  std_logic;
    BA3   : in  std_logic;
    BA4   : in  std_logic;
    BA5   : in  std_logic;
    BA6   : in  std_logic;
    BA7   : in  std_logic;
    BA8   : in  std_logic;
    BA9   : in  std_logic;
    BA10  : in  std_logic;
    BA11  : in  std_logic;
    BA12  : in  std_logic;
    BA13  : in  std_logic;
    BA14  : in  std_logic;
    BA15  : in  std_logic;
    BA16  : in  std_logic;

    BCS   : in  std_logic;
    BWE   : in  std_logic;
    BR    : in  std_logic
);
end NX_RAM_U_BOX;
--#}}}}
-- =================================================================================================
--   NX_DSP_U definition                                                                2020/07/27
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DSP_U is
    generic (
        std_mode    : string                  := "";                             -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
        raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
        raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
        raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
        raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
    );
    port (
        A1    : in std_logic;
        A2    : in std_logic;
        A3    : in std_logic;
        A4    : in std_logic;
        A5    : in std_logic;
        A6    : in std_logic;
        A7    : in std_logic;
        A8    : in std_logic;
        A9    : in std_logic;
        A10   : in std_logic;
        A11   : in std_logic;
        A12   : in std_logic;
        A13   : in std_logic;
        A14   : in std_logic;
        A15   : in std_logic;
        A16   : in std_logic;
        A17   : in std_logic;
        A18   : in std_logic;
        A19   : in std_logic;
        A20   : in std_logic;
        A21   : in std_logic;
        A22   : in std_logic;
        A23   : in std_logic;
        A24   : in std_logic;

        B1    : in std_logic;
        B2    : in std_logic;
        B3    : in std_logic;
        B4    : in std_logic;
        B5    : in std_logic;
        B6    : in std_logic;
        B7    : in std_logic;
        B8    : in std_logic;
        B9    : in std_logic;
        B10   : in std_logic;
        B11   : in std_logic;
        B12   : in std_logic;
        B13   : in std_logic;
        B14   : in std_logic;
        B15   : in std_logic;
        B16   : in std_logic;
        B17   : in std_logic;
        B18   : in std_logic;

        C1    : in std_logic;
        C2    : in std_logic;
        C3    : in std_logic;
        C4    : in std_logic;
        C5    : in std_logic;
        C6    : in std_logic;
        C7    : in std_logic;
        C8    : in std_logic;
        C9    : in std_logic;
        C10   : in std_logic;
        C11   : in std_logic;
        C12   : in std_logic;
        C13   : in std_logic;
        C14   : in std_logic;
        C15   : in std_logic;
        C16   : in std_logic;
        C17   : in std_logic;
        C18   : in std_logic;
        C19   : in std_logic;
        C20   : in std_logic;
        C21   : in std_logic;
        C22   : in std_logic;
        C23   : in std_logic;
        C24   : in std_logic;
        C25   : in std_logic;
        C26   : in std_logic;
        C27   : in std_logic;
        C28   : in std_logic;
        C29   : in std_logic;
        C30   : in std_logic;
        C31   : in std_logic;
        C32   : in std_logic;
        C33   : in std_logic;
        C34   : in std_logic;
        C35   : in std_logic;
        C36   : in std_logic;

        CAI1  : in std_logic;
        CAI2  : in std_logic;
        CAI3  : in std_logic;
        CAI4  : in std_logic;
        CAI5  : in std_logic;
        CAI6  : in std_logic;
        CAI7  : in std_logic;
        CAI8  : in std_logic;
        CAI9  : in std_logic;
        CAI10 : in std_logic;
        CAI11 : in std_logic;
        CAI12 : in std_logic;
        CAI13 : in std_logic;
        CAI14 : in std_logic;
        CAI15 : in std_logic;
        CAI16 : in std_logic;
        CAI17 : in std_logic;
        CAI18 : in std_logic;
        CAI19 : in std_logic;
        CAI20 : in std_logic;
        CAI21 : in std_logic;
        CAI22 : in std_logic;
        CAI23 : in std_logic;
        CAI24 : in std_logic;

        CAO1  : out std_logic;
        CAO2  : out std_logic;
        CAO3  : out std_logic;
        CAO4  : out std_logic;
        CAO5  : out std_logic;
        CAO6  : out std_logic;
        CAO7  : out std_logic;
        CAO8  : out std_logic;
        CAO9  : out std_logic;
        CAO10 : out std_logic;
        CAO11 : out std_logic;
        CAO12 : out std_logic;
        CAO13 : out std_logic;
        CAO14 : out std_logic;
        CAO15 : out std_logic;
        CAO16 : out std_logic;
        CAO17 : out std_logic;
        CAO18 : out std_logic;
        CAO19 : out std_logic;
        CAO20 : out std_logic;
        CAO21 : out std_logic;
        CAO22 : out std_logic;
        CAO23 : out std_logic;
        CAO24 : out std_logic;

        CBI1  : in std_logic;
        CBI2  : in std_logic;
        CBI3  : in std_logic;
        CBI4  : in std_logic;
        CBI5  : in std_logic;
        CBI6  : in std_logic;
        CBI7  : in std_logic;
        CBI8  : in std_logic;
        CBI9  : in std_logic;
        CBI10 : in std_logic;
        CBI11 : in std_logic;
        CBI12 : in std_logic;
        CBI13 : in std_logic;
        CBI14 : in std_logic;
        CBI15 : in std_logic;
        CBI16 : in std_logic;
        CBI17 : in std_logic;
        CBI18 : in std_logic;

        CBO1  : out std_logic;
        CBO2  : out std_logic;
        CBO3  : out std_logic;
        CBO4  : out std_logic;
        CBO5  : out std_logic;
        CBO6  : out std_logic;
        CBO7  : out std_logic;
        CBO8  : out std_logic;
        CBO9  : out std_logic;
        CBO10 : out std_logic;
        CBO11 : out std_logic;
        CBO12 : out std_logic;
        CBO13 : out std_logic;
        CBO14 : out std_logic;
        CBO15 : out std_logic;
        CBO16 : out std_logic;
        CBO17 : out std_logic;
        CBO18 : out std_logic;

        CCI   : in std_logic;
        CCO   : out std_logic;
        CI    : in std_logic;
        CK    : in std_logic;
        CO43  : out std_logic;
        CO57  : out std_logic;
        RESERVED : out std_logic;

        CZI1  : in std_logic;
        CZI2  : in std_logic;
        CZI3  : in std_logic;
        CZI4  : in std_logic;
        CZI5  : in std_logic;
        CZI6  : in std_logic;
        CZI7  : in std_logic;
        CZI8  : in std_logic;
        CZI9  : in std_logic;
        CZI10 : in std_logic;
        CZI11 : in std_logic;
        CZI12 : in std_logic;
        CZI13 : in std_logic;
        CZI14 : in std_logic;
        CZI15 : in std_logic;
        CZI16 : in std_logic;
        CZI17 : in std_logic;
        CZI18 : in std_logic;
        CZI19 : in std_logic;
        CZI20 : in std_logic;
        CZI21 : in std_logic;
        CZI22 : in std_logic;
        CZI23 : in std_logic;
        CZI24 : in std_logic;
        CZI25 : in std_logic;
        CZI26 : in std_logic;
        CZI27 : in std_logic;
        CZI28 : in std_logic;
        CZI29 : in std_logic;
        CZI30 : in std_logic;
        CZI31 : in std_logic;
        CZI32 : in std_logic;
        CZI33 : in std_logic;
        CZI34 : in std_logic;
        CZI35 : in std_logic;
        CZI36 : in std_logic;
        CZI37 : in std_logic;
        CZI38 : in std_logic;
        CZI39 : in std_logic;
        CZI40 : in std_logic;
        CZI41 : in std_logic;
        CZI42 : in std_logic;
        CZI43 : in std_logic;
        CZI44 : in std_logic;
        CZI45 : in std_logic;
        CZI46 : in std_logic;
        CZI47 : in std_logic;
        CZI48 : in std_logic;
        CZI49 : in std_logic;
        CZI50 : in std_logic;
        CZI51 : in std_logic;
        CZI52 : in std_logic;
        CZI53 : in std_logic;
        CZI54 : in std_logic;
        CZI55 : in std_logic;
        CZI56 : in std_logic;

        CZO1  : out std_logic;
        CZO2  : out std_logic;
        CZO3  : out std_logic;
        CZO4  : out std_logic;
        CZO5  : out std_logic;
        CZO6  : out std_logic;
        CZO7  : out std_logic;
        CZO8  : out std_logic;
        CZO9  : out std_logic;
        CZO10 : out std_logic;
        CZO11 : out std_logic;
        CZO12 : out std_logic;
        CZO13 : out std_logic;
        CZO14 : out std_logic;
        CZO15 : out std_logic;
        CZO16 : out std_logic;
        CZO17 : out std_logic;
        CZO18 : out std_logic;
        CZO19 : out std_logic;
        CZO20 : out std_logic;
        CZO21 : out std_logic;
        CZO22 : out std_logic;
        CZO23 : out std_logic;
        CZO24 : out std_logic;
        CZO25 : out std_logic;
        CZO26 : out std_logic;
        CZO27 : out std_logic;
        CZO28 : out std_logic;
        CZO29 : out std_logic;
        CZO30 : out std_logic;
        CZO31 : out std_logic;
        CZO32 : out std_logic;
        CZO33 : out std_logic;
        CZO34 : out std_logic;
        CZO35 : out std_logic;
        CZO36 : out std_logic;
        CZO37 : out std_logic;
        CZO38 : out std_logic;
        CZO39 : out std_logic;
        CZO40 : out std_logic;
        CZO41 : out std_logic;
        CZO42 : out std_logic;
        CZO43 : out std_logic;
        CZO44 : out std_logic;
        CZO45 : out std_logic;
        CZO46 : out std_logic;
        CZO47 : out std_logic;
        CZO48 : out std_logic;
        CZO49 : out std_logic;
        CZO50 : out std_logic;
        CZO51 : out std_logic;
        CZO52 : out std_logic;
        CZO53 : out std_logic;
        CZO54 : out std_logic;
        CZO55 : out std_logic;
        CZO56 : out std_logic;

        D1    : in std_logic;
        D2    : in std_logic;
        D3    : in std_logic;
        D4    : in std_logic;
        D5    : in std_logic;
        D6    : in std_logic;
        D7    : in std_logic;
        D8    : in std_logic;
        D9    : in std_logic;
        D10   : in std_logic;
        D11   : in std_logic;
        D12   : in std_logic;
        D13   : in std_logic;
        D14   : in std_logic;
        D15   : in std_logic;
        D16   : in std_logic;
        D17   : in std_logic;
        D18   : in std_logic;

        OVF   : out std_logic;
        R     : in std_logic;
        RZ    : in std_logic;
        WE    : in std_logic;
        WEZ   : in std_logic;

        Z1    : out std_logic;
        Z2    : out std_logic;
        Z3    : out std_logic;
        Z4    : out std_logic;
        Z5    : out std_logic;
        Z6    : out std_logic;
        Z7    : out std_logic;
        Z8    : out std_logic;
        Z9    : out std_logic;
        Z10   : out std_logic;
        Z11   : out std_logic;
        Z12   : out std_logic;
        Z13   : out std_logic;
        Z14   : out std_logic;
        Z15   : out std_logic;
        Z16   : out std_logic;
        Z17   : out std_logic;
        Z18   : out std_logic;
        Z19   : out std_logic;
        Z20   : out std_logic;
        Z21   : out std_logic;
        Z22   : out std_logic;
        Z23   : out std_logic;
        Z24   : out std_logic;
        Z25   : out std_logic;
        Z26   : out std_logic;
        Z27   : out std_logic;
        Z28   : out std_logic;
        Z29   : out std_logic;
        Z30   : out std_logic;
        Z31   : out std_logic;
        Z32   : out std_logic;
        Z33   : out std_logic;
        Z34   : out std_logic;
        Z35   : out std_logic;
        Z36   : out std_logic;
        Z37   : out std_logic;
        Z38   : out std_logic;
        Z39   : out std_logic;
        Z40   : out std_logic;
        Z41   : out std_logic;
        Z42   : out std_logic;
        Z43   : out std_logic;
        Z44   : out std_logic;
        Z45   : out std_logic;
        Z46   : out std_logic;
        Z47   : out std_logic;
        Z48   : out std_logic;
        Z49   : out std_logic;
        Z50   : out std_logic;
        Z51   : out std_logic;
        Z52   : out std_logic;
        Z53   : out std_logic;
        Z54   : out std_logic;
        Z55   : out std_logic;
        Z56   : out std_logic
    );
end NX_DSP_U;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_U_WRAP definition                                                           2020/07/27
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NX_DSP_U_WRAP is
    generic (
        std_mode    : string                  := "";
        raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
        raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
        raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
        raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
    );
    port (
        A    : in std_logic_vector(23 downto 0);
        B    : in std_logic_vector(17 downto 0);
        C    : in std_logic_vector(35 downto 0);

        CAI  : in std_logic_vector(23 downto 0);
        CAO  : out std_logic_vector(23 downto 0);
        CBI  : in std_logic_vector(17 downto 0);
        CBO  : out std_logic_vector(17 downto 0);

        CCI  : in std_logic;
        CCO  : out std_logic;
        CI   : in std_logic;
        CK   : in std_logic;
        CO43 : out std_logic;
        CO57 : out std_logic;

        CZI  : in std_logic_vector(55 downto 0);
        CZO  : out std_logic_vector(55 downto 0);

        D    : in std_logic_vector(17 downto 0);

        OVF  : out std_logic;
        R    : in std_logic;
        RZ   : in std_logic;
        WE   : in std_logic;
        WEZ  : in std_logic;

        Z    : out std_logic_vector(55 downto 0)
    );
end NX_DSP_U_WRAP;

-- architecture NX_ARCH of NX_DSP_U_WRAP#{{{#
architecture NX_ARCH of NX_DSP_U_WRAP is
    attribute NX_TYPE             : string;
    attribute NX_TYPE of NX_ARCH : architecture is "WRAPPER";

    component NX_DSP_U
        generic (
            std_mode    : string                  := "";
            raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
            raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
            raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
            raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
        );
        port (
            A1    : in std_logic := '0';
            A2    : in std_logic := '0';
            A3    : in std_logic := '0';
            A4    : in std_logic := '0';
            A5    : in std_logic := '0';
            A6    : in std_logic := '0';
            A7    : in std_logic := '0';
            A8    : in std_logic := '0';
            A9    : in std_logic := '0';
            A10   : in std_logic := '0';
            A11   : in std_logic := '0';
            A12   : in std_logic := '0';
            A13   : in std_logic := '0';
            A14   : in std_logic := '0';
            A15   : in std_logic := '0';
            A16   : in std_logic := '0';
            A17   : in std_logic := '0';
            A18   : in std_logic := '0';
            A19   : in std_logic := '0';
            A20   : in std_logic := '0';
            A21   : in std_logic := '0';
            A22   : in std_logic := '0';
            A23   : in std_logic := '0';
            A24   : in std_logic := '0';

            B1    : in std_logic := '0';
            B2    : in std_logic := '0';
            B3    : in std_logic := '0';
            B4    : in std_logic := '0';
            B5    : in std_logic := '0';
            B6    : in std_logic := '0';
            B7    : in std_logic := '0';
            B8    : in std_logic := '0';
            B9    : in std_logic := '0';
            B10   : in std_logic := '0';
            B11   : in std_logic := '0';
            B12   : in std_logic := '0';
            B13   : in std_logic := '0';
            B14   : in std_logic := '0';
            B15   : in std_logic := '0';
            B16   : in std_logic := '0';
            B17   : in std_logic := '0';
            B18   : in std_logic := '0';

            C1    : in std_logic := '0';
            C2    : in std_logic := '0';
            C3    : in std_logic := '0';
            C4    : in std_logic := '0';
            C5    : in std_logic := '0';
            C6    : in std_logic := '0';
            C7    : in std_logic := '0';
            C8    : in std_logic := '0';
            C9    : in std_logic := '0';
            C10   : in std_logic := '0';
            C11   : in std_logic := '0';
            C12   : in std_logic := '0';
            C13   : in std_logic := '0';
            C14   : in std_logic := '0';
            C15   : in std_logic := '0';
            C16   : in std_logic := '0';
            C17   : in std_logic := '0';
            C18   : in std_logic := '0';
            C19   : in std_logic := '0';
            C20   : in std_logic := '0';
            C21   : in std_logic := '0';
            C22   : in std_logic := '0';
            C23   : in std_logic := '0';
            C24   : in std_logic := '0';
            C25   : in std_logic := '0';
            C26   : in std_logic := '0';
            C27   : in std_logic := '0';
            C28   : in std_logic := '0';
            C29   : in std_logic := '0';
            C30   : in std_logic := '0';
            C31   : in std_logic := '0';
            C32   : in std_logic := '0';
            C33   : in std_logic := '0';
            C34   : in std_logic := '0';
            C35   : in std_logic := '0';
            C36   : in std_logic := '0';

            CAI1  : in std_logic := '0';
            CAI2  : in std_logic := '0';
            CAI3  : in std_logic := '0';
            CAI4  : in std_logic := '0';
            CAI5  : in std_logic := '0';
            CAI6  : in std_logic := '0';
            CAI7  : in std_logic := '0';
            CAI8  : in std_logic := '0';
            CAI9  : in std_logic := '0';
            CAI10 : in std_logic := '0';
            CAI11 : in std_logic := '0';
            CAI12 : in std_logic := '0';
            CAI13 : in std_logic := '0';
            CAI14 : in std_logic := '0';
            CAI15 : in std_logic := '0';
            CAI16 : in std_logic := '0';
            CAI17 : in std_logic := '0';
            CAI18 : in std_logic := '0';
            CAI19 : in std_logic := '0';
            CAI20 : in std_logic := '0';
            CAI21 : in std_logic := '0';
            CAI22 : in std_logic := '0';
            CAI23 : in std_logic := '0';
            CAI24 : in std_logic := '0';

            CAO1  : out std_logic := '0';
            CAO2  : out std_logic := '0';
            CAO3  : out std_logic := '0';
            CAO4  : out std_logic := '0';
            CAO5  : out std_logic := '0';
            CAO6  : out std_logic := '0';
            CAO7  : out std_logic := '0';
            CAO8  : out std_logic := '0';
            CAO9  : out std_logic := '0';
            CAO10 : out std_logic := '0';
            CAO11 : out std_logic := '0';
            CAO12 : out std_logic := '0';
            CAO13 : out std_logic := '0';
            CAO14 : out std_logic := '0';
            CAO15 : out std_logic := '0';
            CAO16 : out std_logic := '0';
            CAO17 : out std_logic := '0';
            CAO18 : out std_logic := '0';
            CAO19 : out std_logic := '0';
            CAO20 : out std_logic := '0';
            CAO21 : out std_logic := '0';
            CAO22 : out std_logic := '0';
            CAO23 : out std_logic := '0';
            CAO24 : out std_logic := '0';

            CBI1  : in std_logic := '0';
            CBI2  : in std_logic := '0';
            CBI3  : in std_logic := '0';
            CBI4  : in std_logic := '0';
            CBI5  : in std_logic := '0';
            CBI6  : in std_logic := '0';
            CBI7  : in std_logic := '0';
            CBI8  : in std_logic := '0';
            CBI9  : in std_logic := '0';
            CBI10 : in std_logic := '0';
            CBI11 : in std_logic := '0';
            CBI12 : in std_logic := '0';
            CBI13 : in std_logic := '0';
            CBI14 : in std_logic := '0';
            CBI15 : in std_logic := '0';
            CBI16 : in std_logic := '0';
            CBI17 : in std_logic := '0';
            CBI18 : in std_logic := '0';

            CBO1  : out std_logic := '0';
            CBO2  : out std_logic := '0';
            CBO3  : out std_logic := '0';
            CBO4  : out std_logic := '0';
            CBO5  : out std_logic := '0';
            CBO6  : out std_logic := '0';
            CBO7  : out std_logic := '0';
            CBO8  : out std_logic := '0';
            CBO9  : out std_logic := '0';
            CBO10 : out std_logic := '0';
            CBO11 : out std_logic := '0';
            CBO12 : out std_logic := '0';
            CBO13 : out std_logic := '0';
            CBO14 : out std_logic := '0';
            CBO15 : out std_logic := '0';
            CBO16 : out std_logic := '0';
            CBO17 : out std_logic := '0';
            CBO18 : out std_logic := '0';

            CCI   : in std_logic := '0';
            CCO   : out std_logic := '0';
            CI    : in std_logic := '0';
            CK    : in std_logic := '0';
            CO43  : out std_logic := '0';
            CO57  : out std_logic := '0';
            RESERVED: out std_logic := '0';

            CZI1  : in std_logic := '0';
            CZI2  : in std_logic := '0';
            CZI3  : in std_logic := '0';
            CZI4  : in std_logic := '0';
            CZI5  : in std_logic := '0';
            CZI6  : in std_logic := '0';
            CZI7  : in std_logic := '0';
            CZI8  : in std_logic := '0';
            CZI9  : in std_logic := '0';
            CZI10 : in std_logic := '0';
            CZI11 : in std_logic := '0';
            CZI12 : in std_logic := '0';
            CZI13 : in std_logic := '0';
            CZI14 : in std_logic := '0';
            CZI15 : in std_logic := '0';
            CZI16 : in std_logic := '0';
            CZI17 : in std_logic := '0';
            CZI18 : in std_logic := '0';
            CZI19 : in std_logic := '0';
            CZI20 : in std_logic := '0';
            CZI21 : in std_logic := '0';
            CZI22 : in std_logic := '0';
            CZI23 : in std_logic := '0';
            CZI24 : in std_logic := '0';
            CZI25 : in std_logic := '0';
            CZI26 : in std_logic := '0';
            CZI27 : in std_logic := '0';
            CZI28 : in std_logic := '0';
            CZI29 : in std_logic := '0';
            CZI30 : in std_logic := '0';
            CZI31 : in std_logic := '0';
            CZI32 : in std_logic := '0';
            CZI33 : in std_logic := '0';
            CZI34 : in std_logic := '0';
            CZI35 : in std_logic := '0';
            CZI36 : in std_logic := '0';
            CZI37 : in std_logic := '0';
            CZI38 : in std_logic := '0';
            CZI39 : in std_logic := '0';
            CZI40 : in std_logic := '0';
            CZI41 : in std_logic := '0';
            CZI42 : in std_logic := '0';
            CZI43 : in std_logic := '0';
            CZI44 : in std_logic := '0';
            CZI45 : in std_logic := '0';
            CZI46 : in std_logic := '0';
            CZI47 : in std_logic := '0';
            CZI48 : in std_logic := '0';
            CZI49 : in std_logic := '0';
            CZI50 : in std_logic := '0';
            CZI51 : in std_logic := '0';
            CZI52 : in std_logic := '0';
            CZI53 : in std_logic := '0';
            CZI54 : in std_logic := '0';
            CZI55 : in std_logic := '0';
            CZI56 : in std_logic := '0';

            CZO1  : out std_logic := '0';
            CZO2  : out std_logic := '0';
            CZO3  : out std_logic := '0';
            CZO4  : out std_logic := '0';
            CZO5  : out std_logic := '0';
            CZO6  : out std_logic := '0';
            CZO7  : out std_logic := '0';
            CZO8  : out std_logic := '0';
            CZO9  : out std_logic := '0';
            CZO10 : out std_logic := '0';
            CZO11 : out std_logic := '0';
            CZO12 : out std_logic := '0';
            CZO13 : out std_logic := '0';
            CZO14 : out std_logic := '0';
            CZO15 : out std_logic := '0';
            CZO16 : out std_logic := '0';
            CZO17 : out std_logic := '0';
            CZO18 : out std_logic := '0';
            CZO19 : out std_logic := '0';
            CZO20 : out std_logic := '0';
            CZO21 : out std_logic := '0';
            CZO22 : out std_logic := '0';
            CZO23 : out std_logic := '0';
            CZO24 : out std_logic := '0';
            CZO25 : out std_logic := '0';
            CZO26 : out std_logic := '0';
            CZO27 : out std_logic := '0';
            CZO28 : out std_logic := '0';
            CZO29 : out std_logic := '0';
            CZO30 : out std_logic := '0';
            CZO31 : out std_logic := '0';
            CZO32 : out std_logic := '0';
            CZO33 : out std_logic := '0';
            CZO34 : out std_logic := '0';
            CZO35 : out std_logic := '0';
            CZO36 : out std_logic := '0';
            CZO37 : out std_logic := '0';
            CZO38 : out std_logic := '0';
            CZO39 : out std_logic := '0';
            CZO40 : out std_logic := '0';
            CZO41 : out std_logic := '0';
            CZO42 : out std_logic := '0';
            CZO43 : out std_logic := '0';
            CZO44 : out std_logic := '0';
            CZO45 : out std_logic := '0';
            CZO46 : out std_logic := '0';
            CZO47 : out std_logic := '0';
            CZO48 : out std_logic := '0';
            CZO49 : out std_logic := '0';
            CZO50 : out std_logic := '0';
            CZO51 : out std_logic := '0';
            CZO52 : out std_logic := '0';
            CZO53 : out std_logic := '0';
            CZO54 : out std_logic := '0';
            CZO55 : out std_logic := '0';
            CZO56 : out std_logic := '0';

            D1    : in std_logic := '0';
            D2    : in std_logic := '0';
            D3    : in std_logic := '0';
            D4    : in std_logic := '0';
            D5    : in std_logic := '0';
            D6    : in std_logic := '0';
            D7    : in std_logic := '0';
            D8    : in std_logic := '0';
            D9    : in std_logic := '0';
            D10   : in std_logic := '0';
            D11   : in std_logic := '0';
            D12   : in std_logic := '0';
            D13   : in std_logic := '0';
            D14   : in std_logic := '0';
            D15   : in std_logic := '0';
            D16   : in std_logic := '0';
            D17   : in std_logic := '0';
            D18   : in std_logic := '0';

            OVF   : out std_logic := '0';
            R     : in std_logic := '0';
            RZ    : in std_logic := '0';
            WE    : in std_logic := '0';
            WEZ   : in std_logic := '0';

            Z1    : out std_logic := '0';
            Z2    : out std_logic := '0';
            Z3    : out std_logic := '0';
            Z4    : out std_logic := '0';
            Z5    : out std_logic := '0';
            Z6    : out std_logic := '0';
            Z7    : out std_logic := '0';
            Z8    : out std_logic := '0';
            Z9    : out std_logic := '0';
            Z10   : out std_logic := '0';
            Z11   : out std_logic := '0';
            Z12   : out std_logic := '0';
            Z13   : out std_logic := '0';
            Z14   : out std_logic := '0';
            Z15   : out std_logic := '0';
            Z16   : out std_logic := '0';
            Z17   : out std_logic := '0';
            Z18   : out std_logic := '0';
            Z19   : out std_logic := '0';
            Z20   : out std_logic := '0';
            Z21   : out std_logic := '0';
            Z22   : out std_logic := '0';
            Z23   : out std_logic := '0';
            Z24   : out std_logic := '0';
            Z25   : out std_logic := '0';
            Z26   : out std_logic := '0';
            Z27   : out std_logic := '0';
            Z28   : out std_logic := '0';
            Z29   : out std_logic := '0';
            Z30   : out std_logic := '0';
            Z31   : out std_logic := '0';
            Z32   : out std_logic := '0';
            Z33   : out std_logic := '0';
            Z34   : out std_logic := '0';
            Z35   : out std_logic := '0';
            Z36   : out std_logic := '0';
            Z37   : out std_logic := '0';
            Z38   : out std_logic := '0';
            Z39   : out std_logic := '0';
            Z40   : out std_logic := '0';
            Z41   : out std_logic := '0';
            Z42   : out std_logic := '0';
            Z43   : out std_logic := '0';
            Z44   : out std_logic := '0';
            Z45   : out std_logic := '0';
            Z46   : out std_logic := '0';
            Z47   : out std_logic := '0';
            Z48   : out std_logic := '0';
            Z49   : out std_logic := '0';
            Z50   : out std_logic := '0';
            Z51   : out std_logic := '0';
            Z52   : out std_logic := '0';
            Z53   : out std_logic := '0';
            Z54   : out std_logic := '0';
            Z55   : out std_logic := '0';
            Z56   : out std_logic := '0'
        );
    end component;

begin

    dsp : NX_DSP_U generic map(
        std_mode    => std_mode,
        raw_config0 => raw_config0,
        raw_config1 => raw_config1,
        raw_config2 => raw_config2,
        raw_config3 => raw_config3)
    port map(
        A1    => A(0),
        A2    => A(1),
        A3    => A(2),
        A4    => A(3),
        A5    => A(4),
        A6    => A(5),
        A7    => A(6),
        A8    => A(7),
        A9    => A(8),
        A10   => A(9),
        A11   => A(10),
        A12   => A(11),
        A13   => A(12),
        A14   => A(13),
        A15   => A(14),
        A16   => A(15),
        A17   => A(16),
        A18   => A(17),
        A19   => A(18),
        A20   => A(19),
        A21   => A(20),
        A22   => A(21),
        A23   => A(22),
        A24   => A(23),

        B1    => B(0),
        B2    => B(1),
        B3    => B(2),
        B4    => B(3),
        B5    => B(4),
        B6    => B(5),
        B7    => B(6),
        B8    => B(7),
        B9    => B(8),
        B10   => B(9),
        B11   => B(10),
        B12   => B(11),
        B13   => B(12),
        B14   => B(13),
        B15   => B(14),
        B16   => B(15),
        B17   => B(16),
        B18   => B(17),

        C1    => C(0),
        C2    => C(1),
        C3    => C(2),
        C4    => C(3),
        C5    => C(4),
        C6    => C(5),
        C7    => C(6),
        C8    => C(7),
        C9    => C(8),
        C10   => C(9),
        C11   => C(10),
        C12   => C(11),
        C13   => C(12),
        C14   => C(13),
        C15   => C(14),
        C16   => C(15),
        C17   => C(16),
        C18   => C(17),
        C19   => C(18),
        C20   => C(19),
        C21   => C(20),
        C22   => C(21),
        C23   => C(22),
        C24   => C(23),
        C25   => C(24),
        C26   => C(25),
        C27   => C(26),
        C28   => C(27),
        C29   => C(28),
        C30   => C(29),
        C31   => C(30),
        C32   => C(31),
        C33   => C(32),
        C34   => C(33),
        C35   => C(34),
        C36   => C(35),

        CAI1  => CAI(0),
        CAI2  => CAI(1),
        CAI3  => CAI(2),
        CAI4  => CAI(3),
        CAI5  => CAI(4),
        CAI6  => CAI(5),
        CAI7  => CAI(6),
        CAI8  => CAI(7),
        CAI9  => CAI(8),
        CAI10 => CAI(9),
        CAI11 => CAI(10),
        CAI12 => CAI(11),
        CAI13 => CAI(12),
        CAI14 => CAI(13),
        CAI15 => CAI(14),
        CAI16 => CAI(15),
        CAI17 => CAI(16),
        CAI18 => CAI(17),
        CAI19 => CAI(18),
        CAI20 => CAI(19),
        CAI21 => CAI(20),
        CAI22 => CAI(21),
        CAI23 => CAI(22),
        CAI24 => CAI(23),

        CAO1  => CAO(0),
        CAO2  => CAO(1),
        CAO3  => CAO(2),
        CAO4  => CAO(3),
        CAO5  => CAO(4),
        CAO6  => CAO(5),
        CAO7  => CAO(6),
        CAO8  => CAO(7),
        CAO9  => CAO(8),
        CAO10 => CAO(9),
        CAO11 => CAO(10),
        CAO12 => CAO(11),
        CAO13 => CAO(12),
        CAO14 => CAO(13),
        CAO15 => CAO(14),
        CAO16 => CAO(15),
        CAO17 => CAO(16),
        CAO18 => CAO(17),
        CAO19 => CAO(18),
        CAO20 => CAO(19),
        CAO21 => CAO(20),
        CAO22 => CAO(21),
        CAO23 => CAO(22),
        CAO24 => CAO(23),

        CBI1  => CBI(0),
        CBI2  => CBI(1),
        CBI3  => CBI(2),
        CBI4  => CBI(3),
        CBI5  => CBI(4),
        CBI6  => CBI(5),
        CBI7  => CBI(6),
        CBI8  => CBI(7),
        CBI9  => CBI(8),
        CBI10 => CBI(9),
        CBI11 => CBI(10),
        CBI12 => CBI(11),
        CBI13 => CBI(12),
        CBI14 => CBI(13),
        CBI15 => CBI(14),
        CBI16 => CBI(15),
        CBI17 => CBI(16),
        CBI18 => CBI(17),

        CBO1  => CBO(0),
        CBO2  => CBO(1),
        CBO3  => CBO(2),
        CBO4  => CBO(3),
        CBO5  => CBO(4),
        CBO6  => CBO(5),
        CBO7  => CBO(6),
        CBO8  => CBO(7),
        CBO9  => CBO(8),
        CBO10 => CBO(9),
        CBO11 => CBO(10),
        CBO12 => CBO(11),
        CBO13 => CBO(12),
        CBO14 => CBO(13),
        CBO15 => CBO(14),
        CBO16 => CBO(15),
        CBO17 => CBO(16),
        CBO18 => CBO(17),

        CCI   => CCI,
        CCO   => CCO,
        CI    => CI,
        CK    => CK,
        CO43  => CO43,
        CO57  => CO57,
        RESERVED => OPEN,

        CZI1  => CZI(0),
        CZI2  => CZI(1),
        CZI3  => CZI(2),
        CZI4  => CZI(3),
        CZI5  => CZI(4),
        CZI6  => CZI(5),
        CZI7  => CZI(6),
        CZI8  => CZI(7),
        CZI9  => CZI(8),
        CZI10 => CZI(9),
        CZI11 => CZI(10),
        CZI12 => CZI(11),
        CZI13 => CZI(12),
        CZI14 => CZI(13),
        CZI15 => CZI(14),
        CZI16 => CZI(15),
        CZI17 => CZI(16),
        CZI18 => CZI(17),
        CZI19 => CZI(18),
        CZI20 => CZI(19),
        CZI21 => CZI(20),
        CZI22 => CZI(21),
        CZI23 => CZI(22),
        CZI24 => CZI(23),
        CZI25 => CZI(24),
        CZI26 => CZI(25),
        CZI27 => CZI(26),
        CZI28 => CZI(27),
        CZI29 => CZI(28),
        CZI30 => CZI(29),
        CZI31 => CZI(30),
        CZI32 => CZI(31),
        CZI33 => CZI(32),
        CZI34 => CZI(33),
        CZI35 => CZI(34),
        CZI36 => CZI(35),
        CZI37 => CZI(36),
        CZI38 => CZI(37),
        CZI39 => CZI(38),
        CZI40 => CZI(39),
        CZI41 => CZI(40),
        CZI42 => CZI(41),
        CZI43 => CZI(42),
        CZI44 => CZI(43),
        CZI45 => CZI(44),
        CZI46 => CZI(45),
        CZI47 => CZI(46),
        CZI48 => CZI(47),
        CZI49 => CZI(48),
        CZI50 => CZI(49),
        CZI51 => CZI(50),
        CZI52 => CZI(51),
        CZI53 => CZI(52),
        CZI54 => CZI(53),
        CZI55 => CZI(54),
        CZI56 => CZI(55),

        CZO1  => CZO(0),
        CZO2  => CZO(1),
        CZO3  => CZO(2),
        CZO4  => CZO(3),
        CZO5  => CZO(4),
        CZO6  => CZO(5),
        CZO7  => CZO(6),
        CZO8  => CZO(7),
        CZO9  => CZO(8),
        CZO10 => CZO(9),
        CZO11 => CZO(10),
        CZO12 => CZO(11),
        CZO13 => CZO(12),
        CZO14 => CZO(13),
        CZO15 => CZO(14),
        CZO16 => CZO(15),
        CZO17 => CZO(16),
        CZO18 => CZO(17),
        CZO19 => CZO(18),
        CZO20 => CZO(19),
        CZO21 => CZO(20),
        CZO22 => CZO(21),
        CZO23 => CZO(22),
        CZO24 => CZO(23),
        CZO25 => CZO(24),
        CZO26 => CZO(25),
        CZO27 => CZO(26),
        CZO28 => CZO(27),
        CZO29 => CZO(28),
        CZO30 => CZO(29),
        CZO31 => CZO(30),
        CZO32 => CZO(31),
        CZO33 => CZO(32),
        CZO34 => CZO(33),
        CZO35 => CZO(34),
        CZO36 => CZO(35),
        CZO37 => CZO(36),
        CZO38 => CZO(37),
        CZO39 => CZO(38),
        CZO40 => CZO(39),
        CZO41 => CZO(40),
        CZO42 => CZO(41),
        CZO43 => CZO(42),
        CZO44 => CZO(43),
        CZO45 => CZO(44),
        CZO46 => CZO(45),
        CZO47 => CZO(46),
        CZO48 => CZO(47),
        CZO49 => CZO(48),
        CZO50 => CZO(49),
        CZO51 => CZO(50),
        CZO52 => CZO(51),
        CZO53 => CZO(52),
        CZO54 => CZO(53),
        CZO55 => CZO(54),
        CZO56 => CZO(55),

        D1    => D(0),
        D2    => D(1),
        D3    => D(2),
        D4    => D(3),
        D5    => D(4),
        D6    => D(5),
        D7    => D(6),
        D8    => D(7),
        D9    => D(8),
        D10   => D(9),
        D11   => D(10),
        D12   => D(11),
        D13   => D(12),
        D14   => D(13),
        D15   => D(14),
        D16   => D(15),
        D17   => D(16),
        D18   => D(17),

        OVF   => OVF,
        R     => R,
        RZ    => RZ,
        WE    => WE,
        WEZ   => WEZ,

        Z1    => Z(0),
        Z2    => Z(1),
        Z3    => Z(2),
        Z4    => Z(3),
        Z5    => Z(4),
        Z6    => Z(5),
        Z7    => Z(6),
        Z8    => Z(7),
        Z9    => Z(8),
        Z10   => Z(9),
        Z11   => Z(10),
        Z12   => Z(11),
        Z13   => Z(12),
        Z14   => Z(13),
        Z15   => Z(14),
        Z16   => Z(15),
        Z17   => Z(16),
        Z18   => Z(17),
        Z19   => Z(18),
        Z20   => Z(19),
        Z21   => Z(20),
        Z22   => Z(21),
        Z23   => Z(22),
        Z24   => Z(23),
        Z25   => Z(24),
        Z26   => Z(25),
        Z27   => Z(26),
        Z28   => Z(27),
        Z29   => Z(28),
        Z30   => Z(29),
        Z31   => Z(30),
        Z32   => Z(31),
        Z33   => Z(32),
        Z34   => Z(33),
        Z35   => Z(34),
        Z36   => Z(35),
        Z37   => Z(36),
        Z38   => Z(37),
        Z39   => Z(38),
        Z40   => Z(39),
        Z41   => Z(40),
        Z42   => Z(41),
        Z43   => Z(42),
        Z44   => Z(43),
        Z45   => Z(44),
        Z46   => Z(45),
        Z47   => Z(46),
        Z48   => Z(47),
        Z49   => Z(48),
        Z50   => Z(49),
        Z51   => Z(50),
        Z52   => Z(51),
        Z53   => Z(52),
        Z54   => Z(53),
        Z55   => Z(54),
        Z56   => Z(55)
    );

end NX_ARCH;
-- #}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_DSP_U_SPLIT definition                                                          2020/07/27
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_signed.all;

entity NX_DSP_U_SPLIT is
    generic (
        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config0" (cfg_mode). Defines :
        ------------------------------------------------------------------------- 
        SIGNED_MODE        : bit                    := '0';
        INV_WE             : bit                    := '0';
        INV_WEZ            : bit                    := '0';
        INV_RST            : bit                    := '0';
        INV_RSTZ           : bit                    := '0';
        ALU_DYNAMIC_OP     : bit_vector(1 downto 0) := B"00";     -- "00" for Static,
        -- "-1" for Dynamic control from C
        -- "10" for Dynamic control from D
        SATURATION_RANK    : bit_vector(5 downto 0) := B"000000"; -- Weight of useful MSB on Z and CZO result
        --(to define saturation and overflow)
        ENABLE_SATURATION  : bit                    := '0';       -- '0' for Disable,  '1' for Enable
        MUX_CCO            : bit                    := '0';       -- '0' for CC0 = ALU(42), '1' for CCO = ALU(56)
        MUX_Z              : bit                    := '0';       -- Select Z output. '0' for Y, '1' Saturation / ALU
        MUX_CZ             : bit                    := '0';       -- Select MUX_CZ input. '0' for CZI, '1' for CZO
        MUX_Y              : bit                    := '0';       -- Select ALU's Y input. '0' for MULT output, '1' for (B & A)
        MUX_X              : bit_vector(2 downto 0) := B"000";    -- Select MUX_X operation
        -- "000" for c[33:0]&d[41:34],
        -- "001" for C
        -- "010" for MUX_CZ[39:0]&C[15:0]
        -- "011" for MUX_CZ
        -- "100" for MUX_CZ >> 6
        -- "101" for MUX_CZ >> 12
        -- "110" for MUX_CZ >> 17
        -- "111" for MUX_CZ >> 18
        MUX_CCI            : bit                    := '0';       -- Select '1' input of CI mux. '0' for CCI, '1' for CO_feddback
        MUX_CI             : bit                    := '0';       -- Select input carry of ALU. '0' for CI, '1' for CCI/CO_feedback mux
        MUX_P              : bit                    := '0';       -- '1' for PRE_ADDER, '0' for B input
        MUX_B              : bit                    := '0';       -- '0' = B input, '1' = CBI input
        MUX_A              : bit                    := '0';       -- '0' = A input, '1' = CAI input
        PRE_ADDER_OP       : bit                    := '0';       -- '0' = Additon, '1' = Subraction

        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config1" (cfg_pipe_mux)
        -------------------------------------------------------------------------
        PR_WE_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_WEZ_MUX         : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_RST_MUX         : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_RSTZ_MUX        : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_OV_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_CO_MUX          : bit                    := '0';       -- Registered carry out (CO42 & CO56)
        PR_CCO_MUX         : bit                    := '0';       -- Registered cascade carry out
        PR_Z_MUX           : bit                    := '0';       -- Registered output
        PR_CZ_MUX          : bit                    := '0';       -- Registered cascade output
        PR_Y_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_X_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_CI_MUX          : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_MULT_MUX        : bit                    := '0';       -- No pipe reg  -- Register inside MULT
        PR_P_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg (Pre-adder)
        PR_D_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_C_MUX           : bit                    := '0';       -- '0' for No pipe reg, '1' for 1 pipe reg
        PR_B_CASCADE_MUX   : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels for CAO output. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_B_MUX           : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels on B input. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_A_CASCADE_MUX   : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels for CAO output. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        PR_A_MUX           : bit_vector(1 downto 0) := B"00";     -- Number of pipe reg levels on A input. "-0" for 0 level, "01" for 1 level, "11" for 2 levels
        -------------------------------------------------------------------------
        -- Generic declaration to define the "raw_config2" (cfg_pipe_rst)
        -------------------------------------------------------------------------
        ENABLE_PR_OV_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CO_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CCO_RST  : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_Z_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CZ_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_Y_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_X_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_CI_RST   : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_MULT_RST : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_P_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_D_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_C_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_B_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        ENABLE_PR_A_RST    : bit                    := '0';       -- '0' for Disable, '1' for Enable 
        -- PR_CZ_INIT         : bit_vector(5 downto 0) := B"000000"; -- Value of CZ's pipe register on reset

        -------------------------------------------------------------------------
        -- Constants declaration to define the "cfg_pipe_rst" -- raw_config3(6 downto 0)
        -------------------------------------------------------------------------
        ALU_OP             : bit_vector(2 downto 0) := B"000"     -- ALU operation
        -- x+y+c    = "000"
        -- x-y-c    = "001"
        -- x-y+c-1  = "010"
        -- x+y-c+1  = "011"
        -- -x-y-c-1 = "100"
        -- -x+y+c-1 = "101"
        -- -x+y-c   = "110"
        -- -x-y+c-2 = "111"
    );
    port (
        CK   : in std_logic;
        R    : in std_logic;
        RZ   : in std_logic;
        WE   : in std_logic;
        WEZ  : in std_logic;

        CI   : in std_logic; -- cy_i
        A    : in std_logic_vector(23 downto 0);
        B    : in std_logic_vector(17 downto 0);
        C    : in std_logic_vector(35 downto 0);
        D    : in std_logic_vector(17 downto 0);
        CAI  : in std_logic_vector(23 downto 0);
        CBI  : in std_logic_vector(17 downto 0);
        CZI  : in std_logic_vector(55 downto 0);
        CCI  : in std_logic; -- ccy_i

        Z    : out std_logic_vector(55 downto 0);
        CO42 : out std_logic; -- cy42_o
        CO56 : out std_logic; -- cy56_o
        OVF  : out std_logic;
        CAO  : out std_logic_vector(23 downto 0);
        CBO  : out std_logic_vector(17 downto 0);
        CZO  : out std_logic_vector(55 downto 0);
        CCO  : out std_logic -- ccy_o
    );
end NX_DSP_U_SPLIT;

-- architecture NX_RTL of NX_DSP_U_SPLIT#{{{#
architecture NX_RTL of NX_DSP_U_SPLIT is

    ----------------------------------------------------------
    -- Internal signals to be mapped to the NX_DSP_U component
    ----------------------------------------------------------
        signal A1                : std_logic := '0';
        signal A2                : std_logic := '0';
        signal A3                : std_logic := '0';
        signal A4                : std_logic := '0';
        signal A5                : std_logic := '0';
        signal A6                : std_logic := '0';
        signal A7                : std_logic := '0';
        signal A8                : std_logic := '0';
        signal A9                : std_logic := '0';
        signal A10               : std_logic := '0';
        signal A11               : std_logic := '0';
        signal A12               : std_logic := '0';
        signal A13               : std_logic := '0';
        signal A14               : std_logic := '0';
        signal A15               : std_logic := '0';
        signal A16               : std_logic := '0';
        signal A17               : std_logic := '0';
        signal A18               : std_logic := '0';
        signal A19               : std_logic := '0';
        signal A20               : std_logic := '0';
        signal A21               : std_logic := '0';
        signal A22               : std_logic := '0';
        signal A23               : std_logic := '0';
        signal A24               : std_logic := '0';

        signal B1                : std_logic := '0';
        signal B2                : std_logic := '0';
        signal B3                : std_logic := '0';
        signal B4                : std_logic := '0';
        signal B5                : std_logic := '0';
        signal B6                : std_logic := '0';
        signal B7                : std_logic := '0';
        signal B8                : std_logic := '0';
        signal B9                : std_logic := '0';
        signal B10               : std_logic := '0';
        signal B11               : std_logic := '0';
        signal B12               : std_logic := '0';
        signal B13               : std_logic := '0';
        signal B14               : std_logic := '0';
        signal B15               : std_logic := '0';
        signal B16               : std_logic := '0';
        signal B17               : std_logic := '0';
        signal B18               : std_logic := '0';

        signal C1                : std_logic := '0';
        signal C2                : std_logic := '0';
        signal C3                : std_logic := '0';
        signal C4                : std_logic := '0';
        signal C5                : std_logic := '0';
        signal C6                : std_logic := '0';
        signal C7                : std_logic := '0';
        signal C8                : std_logic := '0';
        signal C9                : std_logic := '0';
        signal C10               : std_logic := '0';
        signal C11               : std_logic := '0';
        signal C12               : std_logic := '0';
        signal C13               : std_logic := '0';
        signal C14               : std_logic := '0';
        signal C15               : std_logic := '0';
        signal C16               : std_logic := '0';
        signal C17               : std_logic := '0';
        signal C18               : std_logic := '0';
        signal C19               : std_logic := '0';
        signal C20               : std_logic := '0';
        signal C21               : std_logic := '0';
        signal C22               : std_logic := '0';
        signal C23               : std_logic := '0';
        signal C24               : std_logic := '0';
        signal C25               : std_logic := '0';
        signal C26               : std_logic := '0';
        signal C27               : std_logic := '0';
        signal C28               : std_logic := '0';
        signal C29               : std_logic := '0';
        signal C30               : std_logic := '0';
        signal C31               : std_logic := '0';
        signal C32               : std_logic := '0';
        signal C33               : std_logic := '0';
        signal C34               : std_logic := '0';
        signal C35               : std_logic := '0';
        signal C36               : std_logic := '0';

        signal CAI1              : std_logic := '0';
        signal CAI2              : std_logic := '0';
        signal CAI3              : std_logic := '0';
        signal CAI4              : std_logic := '0';
        signal CAI5              : std_logic := '0';
        signal CAI6              : std_logic := '0';
        signal CAI7              : std_logic := '0';
        signal CAI8              : std_logic := '0';
        signal CAI9              : std_logic := '0';
        signal CAI10             : std_logic := '0';
        signal CAI11             : std_logic := '0';
        signal CAI12             : std_logic := '0';
        signal CAI13             : std_logic := '0';
        signal CAI14             : std_logic := '0';
        signal CAI15             : std_logic := '0';
        signal CAI16             : std_logic := '0';
        signal CAI17             : std_logic := '0';
        signal CAI18             : std_logic := '0';
        signal CAI19             : std_logic := '0';
        signal CAI20             : std_logic := '0';
        signal CAI21             : std_logic := '0';
        signal CAI22             : std_logic := '0';
        signal CAI23             : std_logic := '0';
        signal CAI24             : std_logic := '0';

        signal CAO1              : std_logic := '0';
        signal CAO2              : std_logic := '0';
        signal CAO3              : std_logic := '0';
        signal CAO4              : std_logic := '0';
        signal CAO5              : std_logic := '0';
        signal CAO6              : std_logic := '0';
        signal CAO7              : std_logic := '0';
        signal CAO8              : std_logic := '0';
        signal CAO9              : std_logic := '0';
        signal CAO10             : std_logic := '0';
        signal CAO11             : std_logic := '0';
        signal CAO12             : std_logic := '0';
        signal CAO13             : std_logic := '0';
        signal CAO14             : std_logic := '0';
        signal CAO15             : std_logic := '0';
        signal CAO16             : std_logic := '0';
        signal CAO17             : std_logic := '0';
        signal CAO18             : std_logic := '0';
        signal CAO19             : std_logic := '0';
        signal CAO20             : std_logic := '0';
        signal CAO21             : std_logic := '0';
        signal CAO22             : std_logic := '0';
        signal CAO23             : std_logic := '0';
        signal CAO24             : std_logic := '0';

        signal CBI1              : std_logic := '0';
        signal CBI2              : std_logic := '0';
        signal CBI3              : std_logic := '0';
        signal CBI4              : std_logic := '0';
        signal CBI5              : std_logic := '0';
        signal CBI6              : std_logic := '0';
        signal CBI7              : std_logic := '0';
        signal CBI8              : std_logic := '0';
        signal CBI9              : std_logic := '0';
        signal CBI10             : std_logic := '0';
        signal CBI11             : std_logic := '0';
        signal CBI12             : std_logic := '0';
        signal CBI13             : std_logic := '0';
        signal CBI14             : std_logic := '0';
        signal CBI15             : std_logic := '0';
        signal CBI16             : std_logic := '0';
        signal CBI17             : std_logic := '0';
        signal CBI18             : std_logic := '0';

        signal CBO1              : std_logic := '0';
        signal CBO2              : std_logic := '0';
        signal CBO3              : std_logic := '0';
        signal CBO4              : std_logic := '0';
        signal CBO5              : std_logic := '0';
        signal CBO6              : std_logic := '0';
        signal CBO7              : std_logic := '0';
        signal CBO8              : std_logic := '0';
        signal CBO9              : std_logic := '0';
        signal CBO10             : std_logic := '0';
        signal CBO11             : std_logic := '0';
        signal CBO12             : std_logic := '0';
        signal CBO13             : std_logic := '0';
        signal CBO14             : std_logic := '0';
        signal CBO15             : std_logic := '0';
        signal CBO16             : std_logic := '0';
        signal CBO17             : std_logic := '0';
        signal CBO18             : std_logic := '0';

        signal CO43              : std_logic := '0';
        signal CO57              : std_logic := '0';

        signal CZI1              : std_logic := '0';
        signal CZI2              : std_logic := '0';
        signal CZI3              : std_logic := '0';
        signal CZI4              : std_logic := '0';
        signal CZI5              : std_logic := '0';
        signal CZI6              : std_logic := '0';
        signal CZI7              : std_logic := '0';
        signal CZI8              : std_logic := '0';
        signal CZI9              : std_logic := '0';
        signal CZI10             : std_logic := '0';
        signal CZI11             : std_logic := '0';
        signal CZI12             : std_logic := '0';
        signal CZI13             : std_logic := '0';
        signal CZI14             : std_logic := '0';
        signal CZI15             : std_logic := '0';
        signal CZI16             : std_logic := '0';
        signal CZI17             : std_logic := '0';
        signal CZI18             : std_logic := '0';
        signal CZI19             : std_logic := '0';
        signal CZI20             : std_logic := '0';
        signal CZI21             : std_logic := '0';
        signal CZI22             : std_logic := '0';
        signal CZI23             : std_logic := '0';
        signal CZI24             : std_logic := '0';
        signal CZI25             : std_logic := '0';
        signal CZI26             : std_logic := '0';
        signal CZI27             : std_logic := '0';
        signal CZI28             : std_logic := '0';
        signal CZI29             : std_logic := '0';
        signal CZI30             : std_logic := '0';
        signal CZI31             : std_logic := '0';
        signal CZI32             : std_logic := '0';
        signal CZI33             : std_logic := '0';
        signal CZI34             : std_logic := '0';
        signal CZI35             : std_logic := '0';
        signal CZI36             : std_logic := '0';
        signal CZI37             : std_logic := '0';
        signal CZI38             : std_logic := '0';
        signal CZI39             : std_logic := '0';
        signal CZI40             : std_logic := '0';
        signal CZI41             : std_logic := '0';
        signal CZI42             : std_logic := '0';
        signal CZI43             : std_logic := '0';
        signal CZI44             : std_logic := '0';
        signal CZI45             : std_logic := '0';
        signal CZI46             : std_logic := '0';
        signal CZI47             : std_logic := '0';
        signal CZI48             : std_logic := '0';
        signal CZI49             : std_logic := '0';
        signal CZI50             : std_logic := '0';
        signal CZI51             : std_logic := '0';
        signal CZI52             : std_logic := '0';
        signal CZI53             : std_logic := '0';
        signal CZI54             : std_logic := '0';
        signal CZI55             : std_logic := '0';
        signal CZI56             : std_logic := '0';

        signal CZO1              : std_logic := '0';
        signal CZO2              : std_logic := '0';
        signal CZO3              : std_logic := '0';
        signal CZO4              : std_logic := '0';
        signal CZO5              : std_logic := '0';
        signal CZO6              : std_logic := '0';
        signal CZO7              : std_logic := '0';
        signal CZO8              : std_logic := '0';
        signal CZO9              : std_logic := '0';
        signal CZO10             : std_logic := '0';
        signal CZO11             : std_logic := '0';
        signal CZO12             : std_logic := '0';
        signal CZO13             : std_logic := '0';
        signal CZO14             : std_logic := '0';
        signal CZO15             : std_logic := '0';
        signal CZO16             : std_logic := '0';
        signal CZO17             : std_logic := '0';
        signal CZO18             : std_logic := '0';
        signal CZO19             : std_logic := '0';
        signal CZO20             : std_logic := '0';
        signal CZO21             : std_logic := '0';
        signal CZO22             : std_logic := '0';
        signal CZO23             : std_logic := '0';
        signal CZO24             : std_logic := '0';
        signal CZO25             : std_logic := '0';
        signal CZO26             : std_logic := '0';
        signal CZO27             : std_logic := '0';
        signal CZO28             : std_logic := '0';
        signal CZO29             : std_logic := '0';
        signal CZO30             : std_logic := '0';
        signal CZO31             : std_logic := '0';
        signal CZO32             : std_logic := '0';
        signal CZO33             : std_logic := '0';
        signal CZO34             : std_logic := '0';
        signal CZO35             : std_logic := '0';
        signal CZO36             : std_logic := '0';
        signal CZO37             : std_logic := '0';
        signal CZO38             : std_logic := '0';
        signal CZO39             : std_logic := '0';
        signal CZO40             : std_logic := '0';
        signal CZO41             : std_logic := '0';
        signal CZO42             : std_logic := '0';
        signal CZO43             : std_logic := '0';
        signal CZO44             : std_logic := '0';
        signal CZO45             : std_logic := '0';
        signal CZO46             : std_logic := '0';
        signal CZO47             : std_logic := '0';
        signal CZO48             : std_logic := '0';
        signal CZO49             : std_logic := '0';
        signal CZO50             : std_logic := '0';
        signal CZO51             : std_logic := '0';
        signal CZO52             : std_logic := '0';
        signal CZO53             : std_logic := '0';
        signal CZO54             : std_logic := '0';
        signal CZO55             : std_logic := '0';
        signal CZO56             : std_logic := '0';

        signal D1                : std_logic := '0';
        signal D2                : std_logic := '0';
        signal D3                : std_logic := '0';
        signal D4                : std_logic := '0';
        signal D5                : std_logic := '0';
        signal D6                : std_logic := '0';
        signal D7                : std_logic := '0';
        signal D8                : std_logic := '0';
        signal D9                : std_logic := '0';
        signal D10               : std_logic := '0';
        signal D11               : std_logic := '0';
        signal D12               : std_logic := '0';
        signal D13               : std_logic := '0';
        signal D14               : std_logic := '0';
        signal D15               : std_logic := '0';
        signal D16               : std_logic := '0';
        signal D17               : std_logic := '0';
        signal D18               : std_logic := '0';

        signal Z1                : std_logic := '0';
        signal Z2                : std_logic := '0';
        signal Z3                : std_logic := '0';
        signal Z4                : std_logic := '0';
        signal Z5                : std_logic := '0';
        signal Z6                : std_logic := '0';
        signal Z7                : std_logic := '0';
        signal Z8                : std_logic := '0';
        signal Z9                : std_logic := '0';
        signal Z10               : std_logic := '0';
        signal Z11               : std_logic := '0';
        signal Z12               : std_logic := '0';
        signal Z13               : std_logic := '0';
        signal Z14               : std_logic := '0';
        signal Z15               : std_logic := '0';
        signal Z16               : std_logic := '0';
        signal Z17               : std_logic := '0';
        signal Z18               : std_logic := '0';
        signal Z19               : std_logic := '0';
        signal Z20               : std_logic := '0';
        signal Z21               : std_logic := '0';
        signal Z22               : std_logic := '0';
        signal Z23               : std_logic := '0';
        signal Z24               : std_logic := '0';
        signal Z25               : std_logic := '0';
        signal Z26               : std_logic := '0';
        signal Z27               : std_logic := '0';
        signal Z28               : std_logic := '0';
        signal Z29               : std_logic := '0';
        signal Z30               : std_logic := '0';
        signal Z31               : std_logic := '0';
        signal Z32               : std_logic := '0';
        signal Z33               : std_logic := '0';
        signal Z34               : std_logic := '0';
        signal Z35               : std_logic := '0';
        signal Z36               : std_logic := '0';
        signal Z37               : std_logic := '0';
        signal Z38               : std_logic := '0';
        signal Z39               : std_logic := '0';
        signal Z40               : std_logic := '0';
        signal Z41               : std_logic := '0';
        signal Z42               : std_logic := '0';
        signal Z43               : std_logic := '0';
        signal Z44               : std_logic := '0';
        signal Z45               : std_logic := '0';
        signal Z46               : std_logic := '0';
        signal Z47               : std_logic := '0';
        signal Z48               : std_logic := '0';
        signal Z49               : std_logic := '0';
        signal Z50               : std_logic := '0';
        signal Z51               : std_logic := '0';
        signal Z52               : std_logic := '0';
        signal Z53               : std_logic := '0';
        signal Z54               : std_logic := '0';
        signal Z55               : std_logic := '0';

    constant raw_config0_gen : bit_vector(26 downto 0)
    := INV_WE & INV_WEZ & INV_RST & INV_RSTZ & MUX_CCO & ALU_DYNAMIC_OP & SATURATION_RANK
     & ENABLE_SATURATION & MUX_Z & MUX_CCI & MUX_CI & MUX_Y & MUX_CZ & MUX_X & MUX_P
     & MUX_B & MUX_A & PRE_ADDER_OP & SIGNED_MODE;

    constant raw_config1_gen : bit_vector(23 downto 0)
    := PR_WE_MUX & PR_WEZ_MUX & PR_RST_MUX & PR_RSTZ_MUX & PR_OV_MUX & PR_CO_MUX & PR_CCO_MUX &
    PR_Z_MUX & PR_CZ_MUX & PR_Y_MUX & PR_X_MUX & PR_CI_MUX & PR_MULT_MUX & PR_P_MUX & PR_D_MUX &
    PR_C_MUX & PR_B_CASCADE_MUX & PR_B_MUX & PR_A_CASCADE_MUX & PR_A_MUX;

    constant raw_config2_gen : bit_vector(13 downto 0)
    := ENABLE_PR_OV_RST & ENABLE_PR_CO_RST & ENABLE_PR_CCO_RST & ENABLE_PR_Z_RST &ENABLE_PR_CZ_RST & 
    ENABLE_PR_MULT_RST &ENABLE_PR_Y_RST & ENABLE_PR_X_RST & ENABLE_PR_P_RST & ENABLE_PR_CI_RST & 
    ENABLE_PR_D_RST & ENABLE_PR_C_RST & ENABLE_PR_B_RST & ENABLE_PR_A_RST;

    constant raw_config3_gen : bit_vector(2 downto 0) := ALU_OP;
    ----------------------------------------------------------
    -- NX_DSP_U declaration
    ----------------------------------------------------------
    component NX_DSP_U
        generic (
            std_mode    : string                  := "";                             -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
            raw_config0 : bit_vector(26 downto 0) := B"000000000000000000000000000"; -- Mux
            raw_config1 : bit_vector(23 downto 0) := B"000000000000000000000000";    -- Pipe Mux
            raw_config2 : bit_vector(13 downto 0) := B"00000000000000";              -- Pipe Reset
            raw_config3 : bit_vector(2 downto 0)  := B"000"                          -- ALU operation
        );
        port (
            A1    : in std_logic  := '0';
            A2    : in std_logic  := '0';
            A3    : in std_logic  := '0';
            A4    : in std_logic  := '0';
            A5    : in std_logic  := '0';
            A6    : in std_logic  := '0';
            A7    : in std_logic  := '0';
            A8    : in std_logic  := '0';
            A9    : in std_logic  := '0';
            A10   : in std_logic  := '0';
            A11   : in std_logic  := '0';
            A12   : in std_logic  := '0';
            A13   : in std_logic  := '0';
            A14   : in std_logic  := '0';
            A15   : in std_logic  := '0';
            A16   : in std_logic  := '0';
            A17   : in std_logic  := '0';
            A18   : in std_logic  := '0';
            A19   : in std_logic  := '0';
            A20   : in std_logic  := '0';
            A21   : in std_logic  := '0';
            A22   : in std_logic  := '0';
            A23   : in std_logic  := '0';
            A24   : in std_logic  := '0';

            B1    : in std_logic  := '0';
            B2    : in std_logic  := '0';
            B3    : in std_logic  := '0';
            B4    : in std_logic  := '0';
            B5    : in std_logic  := '0';
            B6    : in std_logic  := '0';
            B7    : in std_logic  := '0';
            B8    : in std_logic  := '0';
            B9    : in std_logic  := '0';
            B10   : in std_logic  := '0';
            B11   : in std_logic  := '0';
            B12   : in std_logic  := '0';
            B13   : in std_logic  := '0';
            B14   : in std_logic  := '0';
            B15   : in std_logic  := '0';
            B16   : in std_logic  := '0';
            B17   : in std_logic  := '0';
            B18   : in std_logic  := '0';

            C1    : in std_logic  := '0';
            C2    : in std_logic  := '0';
            C3    : in std_logic  := '0';
            C4    : in std_logic  := '0';
            C5    : in std_logic  := '0';
            C6    : in std_logic  := '0';
            C7    : in std_logic  := '0';
            C8    : in std_logic  := '0';
            C9    : in std_logic  := '0';
            C10   : in std_logic  := '0';
            C11   : in std_logic  := '0';
            C12   : in std_logic  := '0';
            C13   : in std_logic  := '0';
            C14   : in std_logic  := '0';
            C15   : in std_logic  := '0';
            C16   : in std_logic  := '0';
            C17   : in std_logic  := '0';
            C18   : in std_logic  := '0';
            C19   : in std_logic  := '0';
            C20   : in std_logic  := '0';
            C21   : in std_logic  := '0';
            C22   : in std_logic  := '0';
            C23   : in std_logic  := '0';
            C24   : in std_logic  := '0';
            C25   : in std_logic  := '0';
            C26   : in std_logic  := '0';
            C27   : in std_logic  := '0';
            C28   : in std_logic  := '0';
            C29   : in std_logic  := '0';
            C30   : in std_logic  := '0';
            C31   : in std_logic  := '0';
            C32   : in std_logic  := '0';
            C33   : in std_logic  := '0';
            C34   : in std_logic  := '0';
            C35   : in std_logic  := '0';
            C36   : in std_logic  := '0';

            CAI1  : in std_logic  := '0';
            CAI2  : in std_logic  := '0';
            CAI3  : in std_logic  := '0';
            CAI4  : in std_logic  := '0';
            CAI5  : in std_logic  := '0';
            CAI6  : in std_logic  := '0';
            CAI7  : in std_logic  := '0';
            CAI8  : in std_logic  := '0';
            CAI9  : in std_logic  := '0';
            CAI10 : in std_logic  := '0';
            CAI11 : in std_logic  := '0';
            CAI12 : in std_logic  := '0';
            CAI13 : in std_logic  := '0';
            CAI14 : in std_logic  := '0';
            CAI15 : in std_logic  := '0';
            CAI16 : in std_logic  := '0';
            CAI17 : in std_logic  := '0';
            CAI18 : in std_logic  := '0';
            CAI19 : in std_logic  := '0';
            CAI20 : in std_logic  := '0';
            CAI21 : in std_logic  := '0';
            CAI22 : in std_logic  := '0';
            CAI23 : in std_logic  := '0';
            CAI24 : in std_logic  := '0';

            CAO1  : out std_logic := '0';
            CAO2  : out std_logic := '0';
            CAO3  : out std_logic := '0';
            CAO4  : out std_logic := '0';
            CAO5  : out std_logic := '0';
            CAO6  : out std_logic := '0';
            CAO7  : out std_logic := '0';
            CAO8  : out std_logic := '0';
            CAO9  : out std_logic := '0';
            CAO10 : out std_logic := '0';
            CAO11 : out std_logic := '0';
            CAO12 : out std_logic := '0';
            CAO13 : out std_logic := '0';
            CAO14 : out std_logic := '0';
            CAO15 : out std_logic := '0';
            CAO16 : out std_logic := '0';
            CAO17 : out std_logic := '0';
            CAO18 : out std_logic := '0';
            CAO19 : out std_logic := '0';
            CAO20 : out std_logic := '0';
            CAO21 : out std_logic := '0';
            CAO22 : out std_logic := '0';
            CAO23 : out std_logic := '0';
            CAO24 : out std_logic := '0';

            CBI1  : in std_logic  := '0';
            CBI2  : in std_logic  := '0';
            CBI3  : in std_logic  := '0';
            CBI4  : in std_logic  := '0';
            CBI5  : in std_logic  := '0';
            CBI6  : in std_logic  := '0';
            CBI7  : in std_logic  := '0';
            CBI8  : in std_logic  := '0';
            CBI9  : in std_logic  := '0';
            CBI10 : in std_logic  := '0';
            CBI11 : in std_logic  := '0';
            CBI12 : in std_logic  := '0';
            CBI13 : in std_logic  := '0';
            CBI14 : in std_logic  := '0';
            CBI15 : in std_logic  := '0';
            CBI16 : in std_logic  := '0';
            CBI17 : in std_logic  := '0';
            CBI18 : in std_logic  := '0';

            CBO1  : out std_logic := '0';
            CBO2  : out std_logic := '0';
            CBO3  : out std_logic := '0';
            CBO4  : out std_logic := '0';
            CBO5  : out std_logic := '0';
            CBO6  : out std_logic := '0';
            CBO7  : out std_logic := '0';
            CBO8  : out std_logic := '0';
            CBO9  : out std_logic := '0';
            CBO10 : out std_logic := '0';
            CBO11 : out std_logic := '0';
            CBO12 : out std_logic := '0';
            CBO13 : out std_logic := '0';
            CBO14 : out std_logic := '0';
            CBO15 : out std_logic := '0';
            CBO16 : out std_logic := '0';
            CBO17 : out std_logic := '0';
            CBO18 : out std_logic := '0';

            CCI   : in std_logic  := '0';
            CCO   : out std_logic := '0';
            CI    : in std_logic  := '0';
            CK    : in std_logic  := '0';
            CO43  : out std_logic := '0';
            CO57  : out std_logic := '0';
            RESERVED: out std_logic := '0';

            CZI1  : in std_logic  := '0';
            CZI2  : in std_logic  := '0';
            CZI3  : in std_logic  := '0';
            CZI4  : in std_logic  := '0';
            CZI5  : in std_logic  := '0';
            CZI6  : in std_logic  := '0';
            CZI7  : in std_logic  := '0';
            CZI8  : in std_logic  := '0';
            CZI9  : in std_logic  := '0';
            CZI10 : in std_logic  := '0';
            CZI11 : in std_logic  := '0';
            CZI12 : in std_logic  := '0';
            CZI13 : in std_logic  := '0';
            CZI14 : in std_logic  := '0';
            CZI15 : in std_logic  := '0';
            CZI16 : in std_logic  := '0';
            CZI17 : in std_logic  := '0';
            CZI18 : in std_logic  := '0';
            CZI19 : in std_logic  := '0';
            CZI20 : in std_logic  := '0';
            CZI21 : in std_logic  := '0';
            CZI22 : in std_logic  := '0';
            CZI23 : in std_logic  := '0';
            CZI24 : in std_logic  := '0';
            CZI25 : in std_logic  := '0';
            CZI26 : in std_logic  := '0';
            CZI27 : in std_logic  := '0';
            CZI28 : in std_logic  := '0';
            CZI29 : in std_logic  := '0';
            CZI30 : in std_logic  := '0';
            CZI31 : in std_logic  := '0';
            CZI32 : in std_logic  := '0';
            CZI33 : in std_logic  := '0';
            CZI34 : in std_logic  := '0';
            CZI35 : in std_logic  := '0';
            CZI36 : in std_logic  := '0';
            CZI37 : in std_logic  := '0';
            CZI38 : in std_logic  := '0';
            CZI39 : in std_logic  := '0';
            CZI40 : in std_logic  := '0';
            CZI41 : in std_logic  := '0';
            CZI42 : in std_logic  := '0';
            CZI43 : in std_logic  := '0';
            CZI44 : in std_logic  := '0';
            CZI45 : in std_logic  := '0';
            CZI46 : in std_logic  := '0';
            CZI47 : in std_logic  := '0';
            CZI48 : in std_logic  := '0';
            CZI49 : in std_logic  := '0';
            CZI50 : in std_logic  := '0';
            CZI51 : in std_logic  := '0';
            CZI52 : in std_logic  := '0';
            CZI53 : in std_logic  := '0';
            CZI54 : in std_logic  := '0';
            CZI55 : in std_logic  := '0';
            CZI56 : in std_logic  := '0';

            CZO1  : out std_logic := '0';
            CZO2  : out std_logic := '0';
            CZO3  : out std_logic := '0';
            CZO4  : out std_logic := '0';
            CZO5  : out std_logic := '0';
            CZO6  : out std_logic := '0';
            CZO7  : out std_logic := '0';
            CZO8  : out std_logic := '0';
            CZO9  : out std_logic := '0';
            CZO10 : out std_logic := '0';
            CZO11 : out std_logic := '0';
            CZO12 : out std_logic := '0';
            CZO13 : out std_logic := '0';
            CZO14 : out std_logic := '0';
            CZO15 : out std_logic := '0';
            CZO16 : out std_logic := '0';
            CZO17 : out std_logic := '0';
            CZO18 : out std_logic := '0';
            CZO19 : out std_logic := '0';
            CZO20 : out std_logic := '0';
            CZO21 : out std_logic := '0';
            CZO22 : out std_logic := '0';
            CZO23 : out std_logic := '0';
            CZO24 : out std_logic := '0';
            CZO25 : out std_logic := '0';
            CZO26 : out std_logic := '0';
            CZO27 : out std_logic := '0';
            CZO28 : out std_logic := '0';
            CZO29 : out std_logic := '0';
            CZO30 : out std_logic := '0';
            CZO31 : out std_logic := '0';
            CZO32 : out std_logic := '0';
            CZO33 : out std_logic := '0';
            CZO34 : out std_logic := '0';
            CZO35 : out std_logic := '0';
            CZO36 : out std_logic := '0';
            CZO37 : out std_logic := '0';
            CZO38 : out std_logic := '0';
            CZO39 : out std_logic := '0';
            CZO40 : out std_logic := '0';
            CZO41 : out std_logic := '0';
            CZO42 : out std_logic := '0';
            CZO43 : out std_logic := '0';
            CZO44 : out std_logic := '0';
            CZO45 : out std_logic := '0';
            CZO46 : out std_logic := '0';
            CZO47 : out std_logic := '0';
            CZO48 : out std_logic := '0';
            CZO49 : out std_logic := '0';
            CZO50 : out std_logic := '0';
            CZO51 : out std_logic := '0';
            CZO52 : out std_logic := '0';
            CZO53 : out std_logic := '0';
            CZO54 : out std_logic := '0';
            CZO55 : out std_logic := '0';
            CZO56 : out std_logic := '0';

            D1    : in std_logic  := '0';
            D2    : in std_logic  := '0';
            D3    : in std_logic  := '0';
            D4    : in std_logic  := '0';
            D5    : in std_logic  := '0';
            D6    : in std_logic  := '0';
            D7    : in std_logic  := '0';
            D8    : in std_logic  := '0';
            D9    : in std_logic  := '0';
            D10   : in std_logic  := '0';
            D11   : in std_logic  := '0';
            D12   : in std_logic  := '0';
            D13   : in std_logic  := '0';
            D14   : in std_logic  := '0';
            D15   : in std_logic  := '0';
            D16   : in std_logic  := '0';
            D17   : in std_logic  := '0';
            D18   : in std_logic  := '0';

            OVF   : out std_logic := '0';
            R     : in std_logic  := '0';
            RZ    : in std_logic  := '0';
            WE    : in std_logic  := '0';
            WEZ   : in std_logic  := '0';

            Z1    : out std_logic := '0';
            Z2    : out std_logic := '0';
            Z3    : out std_logic := '0';
            Z4    : out std_logic := '0';
            Z5    : out std_logic := '0';
            Z6    : out std_logic := '0';
            Z7    : out std_logic := '0';
            Z8    : out std_logic := '0';
            Z9    : out std_logic := '0';
            Z10   : out std_logic := '0';
            Z11   : out std_logic := '0';
            Z12   : out std_logic := '0';
            Z13   : out std_logic := '0';
            Z14   : out std_logic := '0';
            Z15   : out std_logic := '0';
            Z16   : out std_logic := '0';
            Z17   : out std_logic := '0';
            Z18   : out std_logic := '0';
            Z19   : out std_logic := '0';
            Z20   : out std_logic := '0';
            Z21   : out std_logic := '0';
            Z22   : out std_logic := '0';
            Z23   : out std_logic := '0';
            Z24   : out std_logic := '0';
            Z25   : out std_logic := '0';
            Z26   : out std_logic := '0';
            Z27   : out std_logic := '0';
            Z28   : out std_logic := '0';
            Z29   : out std_logic := '0';
            Z30   : out std_logic := '0';
            Z31   : out std_logic := '0';
            Z32   : out std_logic := '0';
            Z33   : out std_logic := '0';
            Z34   : out std_logic := '0';
            Z35   : out std_logic := '0';
            Z36   : out std_logic := '0';
            Z37   : out std_logic := '0';
            Z38   : out std_logic := '0';
            Z39   : out std_logic := '0';
            Z40   : out std_logic := '0';
            Z41   : out std_logic := '0';
            Z42   : out std_logic := '0';
            Z43   : out std_logic := '0';
            Z44   : out std_logic := '0';
            Z45   : out std_logic := '0';
            Z46   : out std_logic := '0';
            Z47   : out std_logic := '0';
            Z48   : out std_logic := '0';
            Z49   : out std_logic := '0';
            Z50   : out std_logic := '0';
            Z51   : out std_logic := '0';
            Z52   : out std_logic := '0';
            Z53   : out std_logic := '0';
            Z54   : out std_logic := '0';
            Z55   : out std_logic := '0';
            Z56   : out std_logic := '0'
        );
    end component;

begin

    ----------------------------------------------------------
    -- Instantiation the NX_DSP_U component
    ----------------------------------------------------------
    DSP_INST : NX_DSP_U
    generic map(
        std_mode    => "",              -- standard mode [ADD36, SUB36, SMUL18, UMUL18, ...] empty for raw
        raw_config0 => raw_config0_gen, -- MODE and MUXes
        raw_config1 => raw_config1_gen, -- Pipeline Registers
        raw_config2 => raw_config2_gen, -- Reset Enable for internal registers
        raw_config3 => raw_config3_gen  -- ALU modes
    )
    port map(
        A1    => A(0),
        A2    => A(1),
        A3    => A(2),
        A4    => A(3),
        A5    => A(4),
        A6    => A(5),
        A7    => A(6),
        A8    => A(7),
        A9    => A(8),
        A10   => A(9),
        A11   => A(10),
        A12   => A(11),
        A13   => A(12),
        A14   => A(13),
        A15   => A(14),
        A16   => A(15),
        A17   => A(16),
        A18   => A(17),
        A19   => A(18),
        A20   => A(19),
        A21   => A(20),
        A22   => A(21),
        A23   => A(22),
        A24   => A(23),

        B1    => B(0),
        B2    => B(1),
        B3    => B(2),
        B4    => B(3),
        B5    => B(4),
        B6    => B(5),
        B7    => B(6),
        B8    => B(7),
        B9    => B(8),
        B10   => B(9),
        B11   => B(10),
        B12   => B(11),
        B13   => B(12),
        B14   => B(13),
        B15   => B(14),
        B16   => B(15),
        B17   => B(16),
        B18   => B(17),

        C1    => C(0),
        C2    => C(1),
        C3    => C(2),
        C4    => C(3),
        C5    => C(4),
        C6    => C(5),
        C7    => C(6),
        C8    => C(7),
        C9    => C(8),
        C10   => C(9),
        C11   => C(10),
        C12   => C(11),
        C13   => C(12),
        C14   => C(13),
        C15   => C(14),
        C16   => C(15),
        C17   => C(16),
        C18   => C(17),
        C19   => C(18),
        C20   => C(19),
        C21   => C(20),
        C22   => C(21),
        C23   => C(22),
        C24   => C(23),
        C25   => C(24),
        C26   => C(25),
        C27   => C(26),
        C28   => C(27),
        C29   => C(28),
        C30   => C(29),
        C31   => C(30),
        C32   => C(31),
        C33   => C(32),
        C34   => C(33),
        C35   => C(34),
        C36   => C(35),

        CAI1  => CAI(0),
        CAI2  => CAI(1),
        CAI3  => CAI(2),
        CAI4  => CAI(3),
        CAI5  => CAI(4),
        CAI6  => CAI(5),
        CAI7  => CAI(6),
        CAI8  => CAI(7),
        CAI9  => CAI(8),
        CAI10 => CAI(9),
        CAI11 => CAI(10),
        CAI12 => CAI(11),
        CAI13 => CAI(12),
        CAI14 => CAI(13),
        CAI15 => CAI(14),
        CAI16 => CAI(15),
        CAI17 => CAI(16),
        CAI18 => CAI(17),
        CAI19 => CAI(18),
        CAI20 => CAI(19),
        CAI21 => CAI(20),
        CAI22 => CAI(21),
        CAI23 => CAI(22),
        CAI24 => CAI(23),

        CAO1  => CAO(0),
        CAO2  => CAO(1),
        CAO3  => CAO(2),
        CAO4  => CAO(3),
        CAO5  => CAO(4),
        CAO6  => CAO(5),
        CAO7  => CAO(6),
        CAO8  => CAO(7),
        CAO9  => CAO(8),
        CAO10 => CAO(9),
        CAO11 => CAO(10),
        CAO12 => CAO(11),
        CAO13 => CAO(12),
        CAO14 => CAO(13),
        CAO15 => CAO(14),
        CAO16 => CAO(15),
        CAO17 => CAO(16),
        CAO18 => CAO(17),
        CAO19 => CAO(18),
        CAO20 => CAO(19),
        CAO21 => CAO(20),
        CAO22 => CAO(21),
        CAO23 => CAO(22),
        CAO24 => CAO(23),

        CBI1  => CBI(0),
        CBI2  => CBI(1),
        CBI3  => CBI(2),
        CBI4  => CBI(3),
        CBI5  => CBI(4),
        CBI6  => CBI(5),
        CBI7  => CBI(6),
        CBI8  => CBI(7),
        CBI9  => CBI(8),
        CBI10 => CBI(9),
        CBI11 => CBI(10),
        CBI12 => CBI(11),
        CBI13 => CBI(12),
        CBI14 => CBI(13),
        CBI15 => CBI(14),
        CBI16 => CBI(15),
        CBI17 => CBI(16),
        CBI18 => CBI(17),

        CBO1  => CBO(0),
        CBO2  => CBO(1),
        CBO3  => CBO(2),
        CBO4  => CBO(3),
        CBO5  => CBO(4),
        CBO6  => CBO(5),
        CBO7  => CBO(6),
        CBO8  => CBO(7),
        CBO9  => CBO(8),
        CBO10 => CBO(9),
        CBO11 => CBO(10),
        CBO12 => CBO(11),
        CBO13 => CBO(12),
        CBO14 => CBO(13),
        CBO15 => CBO(14),
        CBO16 => CBO(15),
        CBO17 => CBO(16),
        CBO18 => CBO(17),

        CCI   => CCI,
        CCO   => CCO,
        CI    => CI,
        CK    => CK,
        CO43  => CO42,
        CO57  => CO56,
        RESERVED => OPEN,

        CZI1  => CZI(0),
        CZI2  => CZI(1),
        CZI3  => CZI(2),
        CZI4  => CZI(3),
        CZI5  => CZI(4),
        CZI6  => CZI(5),
        CZI7  => CZI(6),
        CZI8  => CZI(7),
        CZI9  => CZI(8),
        CZI10 => CZI(9),
        CZI11 => CZI(10),
        CZI12 => CZI(11),
        CZI13 => CZI(12),
        CZI14 => CZI(13),
        CZI15 => CZI(14),
        CZI16 => CZI(15),
        CZI17 => CZI(16),
        CZI18 => CZI(17),
        CZI19 => CZI(18),
        CZI20 => CZI(19),
        CZI21 => CZI(20),
        CZI22 => CZI(21),
        CZI23 => CZI(22),
        CZI24 => CZI(23),
        CZI25 => CZI(24),
        CZI26 => CZI(25),
        CZI27 => CZI(26),
        CZI28 => CZI(27),
        CZI29 => CZI(28),
        CZI30 => CZI(29),
        CZI31 => CZI(30),
        CZI32 => CZI(31),
        CZI33 => CZI(32),
        CZI34 => CZI(33),
        CZI35 => CZI(34),
        CZI36 => CZI(35),
        CZI37 => CZI(36),
        CZI38 => CZI(37),
        CZI39 => CZI(38),
        CZI40 => CZI(39),
        CZI41 => CZI(40),
        CZI42 => CZI(41),
        CZI43 => CZI(42),
        CZI44 => CZI(43),
        CZI45 => CZI(44),
        CZI46 => CZI(45),
        CZI47 => CZI(46),
        CZI48 => CZI(47),
        CZI49 => CZI(48),
        CZI50 => CZI(49),
        CZI51 => CZI(50),
        CZI52 => CZI(51),
        CZI53 => CZI(52),
        CZI54 => CZI(53),
        CZI55 => CZI(54),
        CZI56 => CZI(55),

        CZO1  => CZO(0),
        CZO2  => CZO(1),
        CZO3  => CZO(2),
        CZO4  => CZO(3),
        CZO5  => CZO(4),
        CZO6  => CZO(5),
        CZO7  => CZO(6),
        CZO8  => CZO(7),
        CZO9  => CZO(8),
        CZO10 => CZO(9),
        CZO11 => CZO(10),
        CZO12 => CZO(11),
        CZO13 => CZO(12),
        CZO14 => CZO(13),
        CZO15 => CZO(14),
        CZO16 => CZO(15),
        CZO17 => CZO(16),
        CZO18 => CZO(17),
        CZO19 => CZO(18),
        CZO20 => CZO(19),
        CZO21 => CZO(20),
        CZO22 => CZO(21),
        CZO23 => CZO(22),
        CZO24 => CZO(23),
        CZO25 => CZO(24),
        CZO26 => CZO(25),
        CZO27 => CZO(26),
        CZO28 => CZO(27),
        CZO29 => CZO(28),
        CZO30 => CZO(29),
        CZO31 => CZO(30),
        CZO32 => CZO(31),
        CZO33 => CZO(32),
        CZO34 => CZO(33),
        CZO35 => CZO(34),
        CZO36 => CZO(35),
        CZO37 => CZO(36),
        CZO38 => CZO(37),
        CZO39 => CZO(38),
        CZO40 => CZO(39),
        CZO41 => CZO(40),
        CZO42 => CZO(41),
        CZO43 => CZO(42),
        CZO44 => CZO(43),
        CZO45 => CZO(44),
        CZO46 => CZO(45),
        CZO47 => CZO(46),
        CZO48 => CZO(47),
        CZO49 => CZO(48),
        CZO50 => CZO(49),
        CZO51 => CZO(50),
        CZO52 => CZO(51),
        CZO53 => CZO(52),
        CZO54 => CZO(53),
        CZO55 => CZO(54),
        CZO56 => CZO(55),

        D1    => D(0),
        D2    => D(1),
        D3    => D(2),
        D4    => D(3),
        D5    => D(4),
        D6    => D(5),
        D7    => D(6),
        D8    => D(7),
        D9    => D(8),
        D10   => D(9),
        D11   => D(10),
        D12   => D(11),
        D13   => D(12),
        D14   => D(13),
        D15   => D(14),
        D16   => D(15),
        D17   => D(16),
        D18   => D(17),

        OVF   => OVF,
        R     => R,
        RZ    => RZ,
        WE    => WE,

        Z1    => Z(0),
        Z2    => Z(1),
        Z3    => Z(2),
        Z4    => Z(3),
        Z5    => Z(4),
        Z6    => Z(5),
        Z7    => Z(6),
        Z8    => Z(7),
        Z9    => Z(8),
        Z10   => Z(9),
        Z11   => Z(10),
        Z12   => Z(11),
        Z13   => Z(12),
        Z14   => Z(13),
        Z15   => Z(14),
        Z16   => Z(15),
        Z17   => Z(16),
        Z18   => Z(17),
        Z19   => Z(18),
        Z20   => Z(19),
        Z21   => Z(20),
        Z22   => Z(21),
        Z23   => Z(22),
        Z24   => Z(23),
        Z25   => Z(24),
        Z26   => Z(25),
        Z27   => Z(26),
        Z28   => Z(27),
        Z29   => Z(28),
        Z30   => Z(29),
        Z31   => Z(30),
        Z32   => Z(31),
        Z33   => Z(32),
        Z34   => Z(33),
        Z35   => Z(34),
        Z36   => Z(35),
        Z37   => Z(36),
        Z38   => Z(37),
        Z39   => Z(38),
        Z40   => Z(39),
        Z41   => Z(40),
        Z42   => Z(41),
        Z43   => Z(42),
        Z44   => Z(43),
        Z45   => Z(44),
        Z46   => Z(45),
        Z47   => Z(46),
        Z48   => Z(47),
        Z49   => Z(48),
        Z50   => Z(49),
        Z51   => Z(50),
        Z52   => Z(51),
        Z53   => Z(52),
        Z54   => Z(53),
        Z55   => Z(54),
        Z56   => Z(55)
    );

end NX_RTL;
-- #}}}#
-- =================================================================================================
--   NX_FIFO definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_FIFO is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(5 downto 0) := "000000"
);
port (
    RCK   : in  std_logic;
    WCK   : in  std_logic;
    WE    : in  std_logic;
    WEA   : in  std_logic;
    I     : in  std_logic_vector(17 downto 0);
    O     : out std_logic_vector(17 downto 0);
    WRSTI : in  std_logic;
    WAI   : in  std_logic_vector(5 downto 0);
    WAO   : out std_logic_vector(5 downto 0);
    WEQ   : out std_logic;
    RRSTI : in  std_logic;
    RAI   : in  std_logic_vector(5 downto 0);
    RAO   : out std_logic_vector(5 downto 0);
    REQ   : out std_logic
);
end NX_FIFO;

architecture NX_RTL of NX_FIFO is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_FIFO_U
generic (
    mode           : integer := 0;
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK    : in  std_logic;
    WCK    : in  std_logic;
    WE     : in  std_logic;
    WEA    : in  std_logic;
    I1     : in  std_logic;
    I2     : in  std_logic;
    I3     : in  std_logic;
    I4     : in  std_logic;
    I5     : in  std_logic;
    I6     : in  std_logic;
    I7     : in  std_logic;
    I8     : in  std_logic;
    I9     : in  std_logic;
    I10    : in  std_logic;
    I11    : in  std_logic;
    I12    : in  std_logic;
    I13    : in  std_logic;
    I14    : in  std_logic;
    I15    : in  std_logic;
    I16    : in  std_logic;
    I17    : in  std_logic;
    I18    : in  std_logic;
    I19    : in  std_logic;
    I20    : in  std_logic;
    I21    : in  std_logic;
    I22    : in  std_logic;
    I23    : in  std_logic;
    I24    : in  std_logic;
    I25    : in  std_logic;
    I26    : in  std_logic;
    I27    : in  std_logic;
    I28    : in  std_logic;
    I29    : in  std_logic;
    I30    : in  std_logic;
    I31    : in  std_logic;
    I32    : in  std_logic;
    I33    : in  std_logic;
    I34    : in  std_logic;
    I35    : in  std_logic;
    I36    : in  std_logic;
    O1     : out std_logic;
    O2     : out std_logic;
    O3     : out std_logic;
    O4     : out std_logic;
    O5     : out std_logic;
    O6     : out std_logic;
    O7     : out std_logic;
    O8     : out std_logic;
    O9     : out std_logic;
    O10    : out std_logic;
    O11    : out std_logic;
    O12    : out std_logic;
    O13    : out std_logic;
    O14    : out std_logic;
    O15    : out std_logic;
    O16    : out std_logic;
    O17    : out std_logic;
    O18    : out std_logic;
    O19    : out std_logic;
    O20    : out std_logic;
    O21    : out std_logic;
    O22    : out std_logic;
    O23    : out std_logic;
    O24    : out std_logic;
    O25    : out std_logic;
    O26    : out std_logic;
    O27    : out std_logic;
    O28    : out std_logic;
    O29    : out std_logic;
    O30    : out std_logic;
    O31    : out std_logic;
    O32    : out std_logic;
    O33    : out std_logic;
    O34    : out std_logic;
    O35    : out std_logic;
    O36    : out std_logic;
    WRSTI  : in  std_logic;
    WAI1   : in  std_logic;
    WAI2   : in  std_logic;
    WAI3   : in  std_logic;
    WAI4   : in  std_logic;
    WAI5   : in  std_logic;
    WAI6   : in  std_logic;
    WAI7   : in  std_logic;
    WAO1   : out std_logic;
    WAO2   : out std_logic;
    WAO3   : out std_logic;
    WAO4   : out std_logic;
    WAO5   : out std_logic;
    WAO6   : out std_logic;
    WAO7   : out std_logic;
    WEQ1   : out std_logic;
    WEQ2   : out std_logic;
    RRSTI  : in  std_logic;
    RAI1   : in  std_logic;
    RAI2   : in  std_logic;
    RAI3   : in  std_logic;
    RAI4   : in  std_logic;
    RAI5   : in  std_logic;
    RAI6   : in  std_logic;
    RAI7   : in  std_logic;
    RAO1   : out std_logic;
    RAO2   : out std_logic;
    RAO3   : out std_logic;
    RAO4   : out std_logic;
    RAO5   : out std_logic;
    RAO6   : out std_logic;
    RAO7   : out std_logic;
    REQ1   : out std_logic;
    REQ2   : out std_logic
);
end component NX_FIFO_U;

begin

fifo: NX_FIFO_U
generic map (
    mode           => 0, -- 0: DPREG
    wck_edge       => wck_edge,
    rck_edge       => rck_edge,
    use_write_arst => use_write_arst,
    use_read_arst  => use_read_arst
)
port map (
    RCK   => RCK,
    WCK   => WCK,
    WE    => WE,
    WEA   => WEA,
    I1    => I(0),
    I2    => I(1),
    I3    => I(2),
    I4    => I(3),
    I5    => I(4),
    I6    => I(5),
    I7    => I(6),
    I8    => I(7),
    I9    => I(8),
    I10   => I(9),
    I11   => I(10),
    I12   => I(11),
    I13   => I(12),
    I14   => I(13),
    I15   => I(14),
    I16   => I(15),
    I17   => I(16),
    I18   => I(17),
    I19   => '0',
    I20   => '0',
    I21   => '0',
    I22   => '0',
    I23   => '0',
    I24   => '0',
    I25   => '0',
    I26   => '0',
    I27   => '0',
    I28   => '0',
    I29   => '0',
    I30   => '0',
    I31   => '0',
    I32   => '0',
    I33   => '0',
    I34   => '0',
    I35   => '0',
    I36   => '0',
    O1    => O(0),
    O2    => O(1),
    O3    => O(2),
    O4    => O(3),
    O5    => O(4),
    O6    => O(5),
    O7    => O(6),
    O8    => O(7),
    O9    => O(8),
    O10   => O(9),
    O11   => O(10),
    O12   => O(11),
    O13   => O(12),
    O14   => O(13),
    O15   => O(14),
    O16   => O(15),
    O17   => O(16),
    O18   => O(17),
    O19   => OPEN,
    O20   => OPEN,
    O21   => OPEN,
    O22   => OPEN,
    O23   => OPEN,
    O24   => OPEN,
    O25   => OPEN,
    O26   => OPEN,
    O27   => OPEN,
    O28   => OPEN,
    O29   => OPEN,
    O30   => OPEN,
    O31   => OPEN,
    O32   => OPEN,
    O33   => OPEN,
    O34   => OPEN,
    O35   => OPEN,
    O36   => OPEN,
    WRSTI => WRSTI,
    WAI1  => WAI(0),
    WAI2  => WAI(1),
    WAI3  => WAI(2),
    WAI4  => WAI(3),
    WAI5  => WAI(4),
    WAI6  => WAI(5),
    WAI7  => '0',
    WAO1  => WAO(0),
    WAO2  => WAO(1),
    WAO3  => WAO(2),
    WAO4  => WAO(3),
    WAO5  => WAO(4),
    WAO6  => WAO(5),
    WAO7  => OPEN,
    WEQ1  => WEQ,
    WEQ2  => OPEN,
    RRSTI => RRSTI,
    RAI1  => RAI(0),
    RAI2  => RAI(1),
    RAI3  => RAI(2),
    RAI4  => RAI(3),
    RAI5  => RAI(4),
    RAI6  => RAI(5),
    RAI7  => '0',
    RAO1  => RAO(0),
    RAO2  => RAO(1),
    RAO3  => RAO(2),
    RAO4  => RAO(3),
    RAO5  => RAO(4),
    RAO6  => RAO(5),
    RAO7  => OPEN,
    REQ1  => REQ,
    REQ2  => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_XFIFO_64x18 definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XFIFO_64x18 is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK   : in  std_logic;
    WCK   : in  std_logic;
    WE    : in  std_logic;
    WEA   : in  std_logic;
    I     : in  std_logic_vector(17 downto 0);
    O     : out std_logic_vector(17 downto 0);
    WRSTI : in  std_logic;
    WAI   : in  std_logic_vector(6 downto 0);
    WAO   : out std_logic_vector(6 downto 0);
    WEQ   : out std_logic_vector(1 downto 0);
    RRSTI : in  std_logic;
    RAI   : in  std_logic_vector(6 downto 0);
    RAO   : out std_logic_vector(6 downto 0);
    REQ   : out std_logic_vector(1 downto 0)
);
end NX_XFIFO_64x18;

architecture NX_RTL of NX_XFIFO_64x18 is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_FIFO_U
generic (
    mode           : integer := 0;
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK    : in  std_logic;
    WCK    : in  std_logic;
    WE     : in  std_logic;
    WEA    : in  std_logic;
    I1     : in  std_logic;
    I2     : in  std_logic;
    I3     : in  std_logic;
    I4     : in  std_logic;
    I5     : in  std_logic;
    I6     : in  std_logic;
    I7     : in  std_logic;
    I8     : in  std_logic;
    I9     : in  std_logic;
    I10    : in  std_logic;
    I11    : in  std_logic;
    I12    : in  std_logic;
    I13    : in  std_logic;
    I14    : in  std_logic;
    I15    : in  std_logic;
    I16    : in  std_logic;
    I17    : in  std_logic;
    I18    : in  std_logic;
    I19    : in  std_logic;
    I20    : in  std_logic;
    I21    : in  std_logic;
    I22    : in  std_logic;
    I23    : in  std_logic;
    I24    : in  std_logic;
    I25    : in  std_logic;
    I26    : in  std_logic;
    I27    : in  std_logic;
    I28    : in  std_logic;
    I29    : in  std_logic;
    I30    : in  std_logic;
    I31    : in  std_logic;
    I32    : in  std_logic;
    I33    : in  std_logic;
    I34    : in  std_logic;
    I35    : in  std_logic;
    I36    : in  std_logic;
    O1     : out std_logic;
    O2     : out std_logic;
    O3     : out std_logic;
    O4     : out std_logic;
    O5     : out std_logic;
    O6     : out std_logic;
    O7     : out std_logic;
    O8     : out std_logic;
    O9     : out std_logic;
    O10    : out std_logic;
    O11    : out std_logic;
    O12    : out std_logic;
    O13    : out std_logic;
    O14    : out std_logic;
    O15    : out std_logic;
    O16    : out std_logic;
    O17    : out std_logic;
    O18    : out std_logic;
    O19    : out std_logic;
    O20    : out std_logic;
    O21    : out std_logic;
    O22    : out std_logic;
    O23    : out std_logic;
    O24    : out std_logic;
    O25    : out std_logic;
    O26    : out std_logic;
    O27    : out std_logic;
    O28    : out std_logic;
    O29    : out std_logic;
    O30    : out std_logic;
    O31    : out std_logic;
    O32    : out std_logic;
    O33    : out std_logic;
    O34    : out std_logic;
    O35    : out std_logic;
    O36    : out std_logic;
    WRSTI  : in  std_logic;
    WAI1   : in  std_logic;
    WAI2   : in  std_logic;
    WAI3   : in  std_logic;
    WAI4   : in  std_logic;
    WAI5   : in  std_logic;
    WAI6   : in  std_logic;
    WAI7   : in  std_logic;
    WAO1   : out std_logic;
    WAO2   : out std_logic;
    WAO3   : out std_logic;
    WAO4   : out std_logic;
    WAO5   : out std_logic;
    WAO6   : out std_logic;
    WAO7   : out std_logic;
    WEQ1   : out std_logic;
    WEQ2   : out std_logic;
    RRSTI  : in  std_logic;
    RAI1   : in  std_logic;
    RAI2   : in  std_logic;
    RAI3   : in  std_logic;
    RAI4   : in  std_logic;
    RAI5   : in  std_logic;
    RAI6   : in  std_logic;
    RAI7   : in  std_logic;
    RAO1   : out std_logic;
    RAO2   : out std_logic;
    RAO3   : out std_logic;
    RAO4   : out std_logic;
    RAO5   : out std_logic;
    RAO6   : out std_logic;
    RAO7   : out std_logic;
    REQ1   : out std_logic;
    REQ2   : out std_logic
);
end component NX_FIFO_U;

begin

fifo: NX_FIFO_U
generic map (
    mode           => 1, -- 1: XFIFO_64x18
    wck_edge       => wck_edge,
    rck_edge       => rck_edge,
    use_write_arst => use_write_arst,
    use_read_arst  => use_read_arst
)
port map (
    RCK   => RCK,
    WCK   => WCK,
    WE    => WE,
    WEA   => WEA,
    I1    => I(0),
    I2    => I(1),
    I3    => I(2),
    I4    => I(3),
    I5    => I(4),
    I6    => I(5),
    I7    => I(6),
    I8    => I(7),
    I9    => I(8),
    I10   => I(9),
    I11   => I(10),
    I12   => I(11),
    I13   => I(12),
    I14   => I(13),
    I15   => I(14),
    I16   => I(15),
    I17   => I(16),
    I18   => I(17),
    I19   => '0',
    I20   => '0',
    I21   => '0',
    I22   => '0',
    I23   => '0',
    I24   => '0',
    I25   => '0',
    I26   => '0',
    I27   => '0',
    I28   => '0',
    I29   => '0',
    I30   => '0',
    I31   => '0',
    I32   => '0',
    I33   => '0',
    I34   => '0',
    I35   => '0',
    I36   => '0',
    O1    => O(0),
    O2    => O(1),
    O3    => O(2),
    O4    => O(3),
    O5    => O(4),
    O6    => O(5),
    O7    => O(6),
    O8    => O(7),
    O9    => O(8),
    O10   => O(9),
    O11   => O(10),
    O12   => O(11),
    O13   => O(12),
    O14   => O(13),
    O15   => O(14),
    O16   => O(15),
    O17   => O(16),
    O18   => O(17),
    O19   => OPEN,
    O20   => OPEN,
    O21   => OPEN,
    O22   => OPEN,
    O23   => OPEN,
    O24   => OPEN,
    O25   => OPEN,
    O26   => OPEN,
    O27   => OPEN,
    O28   => OPEN,
    O29   => OPEN,
    O30   => OPEN,
    O31   => OPEN,
    O32   => OPEN,
    O33   => OPEN,
    O34   => OPEN,
    O35   => OPEN,
    O36   => OPEN,
    WRSTI => WRSTI,
    WAI1  => WAI(0),
    WAI2  => WAI(1),
    WAI3  => WAI(2),
    WAI4  => WAI(3),
    WAI5  => WAI(4),
    WAI6  => WAI(5),
    WAI7  => WAI(6),
    WAO1  => WAO(0),
    WAO2  => WAO(1),
    WAO3  => WAO(2),
    WAO4  => WAO(3),
    WAO5  => WAO(4),
    WAO6  => WAO(5),
    WAO7  => WAO(6),
    WEQ1  => WEQ(0),
    WEQ2  => WEQ(1),
    RRSTI => RRSTI,
    RAI1  => RAI(0),
    RAI2  => RAI(1),
    RAI3  => RAI(2),
    RAI4  => RAI(3),
    RAI5  => RAI(4),
    RAI6  => RAI(5),
    RAI7  => RAI(6),
    RAO1  => RAO(0),
    RAO2  => RAO(1),
    RAO3  => RAO(2),
    RAO4  => RAO(3),
    RAO5  => RAO(4),
    RAO6  => RAO(5),
    RAO7  => RAO(6),
    REQ1  => REQ(0),
    REQ2  => REQ(1)
);
end NX_RTL;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_XFIFO_32x36 definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XFIFO_32x36 is
generic (
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK   : in  std_logic;
    WCK   : in  std_logic;
    WE    : in  std_logic;
    WEA   : in  std_logic;
    I     : in  std_logic_vector(35 downto 0);
    O     : out std_logic_vector(35 downto 0);
    WRSTI : in  std_logic;
    WAI   : in  std_logic_vector(5 downto 0);
    WAO   : out std_logic_vector(5 downto 0);
    WEQ   : out std_logic;
    RRSTI : in  std_logic;
    RAI   : in  std_logic_vector(5 downto 0);
    RAO   : out std_logic_vector(5 downto 0);
    REQ   : out std_logic
);
end NX_XFIFO_32x36;

architecture NX_RTL of NX_XFIFO_32x36 is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_FIFO_U
generic (
    mode           : integer := 0;
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK    : in  std_logic;
    WCK    : in  std_logic;
    WE     : in  std_logic;
    WEA    : in  std_logic;
    I1     : in  std_logic;
    I2     : in  std_logic;
    I3     : in  std_logic;
    I4     : in  std_logic;
    I5     : in  std_logic;
    I6     : in  std_logic;
    I7     : in  std_logic;
    I8     : in  std_logic;
    I9     : in  std_logic;
    I10    : in  std_logic;
    I11    : in  std_logic;
    I12    : in  std_logic;
    I13    : in  std_logic;
    I14    : in  std_logic;
    I15    : in  std_logic;
    I16    : in  std_logic;
    I17    : in  std_logic;
    I18    : in  std_logic;
    I19    : in  std_logic;
    I20    : in  std_logic;
    I21    : in  std_logic;
    I22    : in  std_logic;
    I23    : in  std_logic;
    I24    : in  std_logic;
    I25    : in  std_logic;
    I26    : in  std_logic;
    I27    : in  std_logic;
    I28    : in  std_logic;
    I29    : in  std_logic;
    I30    : in  std_logic;
    I31    : in  std_logic;
    I32    : in  std_logic;
    I33    : in  std_logic;
    I34    : in  std_logic;
    I35    : in  std_logic;
    I36    : in  std_logic;
    O1     : out std_logic;
    O2     : out std_logic;
    O3     : out std_logic;
    O4     : out std_logic;
    O5     : out std_logic;
    O6     : out std_logic;
    O7     : out std_logic;
    O8     : out std_logic;
    O9     : out std_logic;
    O10    : out std_logic;
    O11    : out std_logic;
    O12    : out std_logic;
    O13    : out std_logic;
    O14    : out std_logic;
    O15    : out std_logic;
    O16    : out std_logic;
    O17    : out std_logic;
    O18    : out std_logic;
    O19    : out std_logic;
    O20    : out std_logic;
    O21    : out std_logic;
    O22    : out std_logic;
    O23    : out std_logic;
    O24    : out std_logic;
    O25    : out std_logic;
    O26    : out std_logic;
    O27    : out std_logic;
    O28    : out std_logic;
    O29    : out std_logic;
    O30    : out std_logic;
    O31    : out std_logic;
    O32    : out std_logic;
    O33    : out std_logic;
    O34    : out std_logic;
    O35    : out std_logic;
    O36    : out std_logic;
    WRSTI  : in  std_logic;
    WAI1   : in  std_logic;
    WAI2   : in  std_logic;
    WAI3   : in  std_logic;
    WAI4   : in  std_logic;
    WAI5   : in  std_logic;
    WAI6   : in  std_logic;
    WAI7   : in  std_logic;
    WAO1   : out std_logic;
    WAO2   : out std_logic;
    WAO3   : out std_logic;
    WAO4   : out std_logic;
    WAO5   : out std_logic;
    WAO6   : out std_logic;
    WAO7   : out std_logic;
    WEQ1   : out std_logic;
    WEQ2   : out std_logic;
    RRSTI  : in  std_logic;
    RAI1   : in  std_logic;
    RAI2   : in  std_logic;
    RAI3   : in  std_logic;
    RAI4   : in  std_logic;
    RAI5   : in  std_logic;
    RAI6   : in  std_logic;
    RAI7   : in  std_logic;
    RAO1   : out std_logic;
    RAO2   : out std_logic;
    RAO3   : out std_logic;
    RAO4   : out std_logic;
    RAO5   : out std_logic;
    RAO6   : out std_logic;
    RAO7   : out std_logic;
    REQ1   : out std_logic;
    REQ2   : out std_logic
);
end component NX_FIFO_U;

begin

fifo: NX_FIFO_U
generic map (
    mode           => 2, -- 2: XFIFO_32x36
    wck_edge       => wck_edge,
    rck_edge       => rck_edge,
    use_write_arst => use_write_arst,
    use_read_arst  => use_read_arst
)
port map (
    RCK   => RCK,
    WCK   => WCK,
    WE    => WE,
    WEA   => WEA,
    I1    => I(0),
    I2    => I(1),
    I3    => I(2),
    I4    => I(3),
    I5    => I(4),
    I6    => I(5),
    I7    => I(6),
    I8    => I(7),
    I9    => I(8),
    I10   => I(9),
    I11   => I(10),
    I12   => I(11),
    I13   => I(12),
    I14   => I(13),
    I15   => I(14),
    I16   => I(15),
    I17   => I(16),
    I18   => I(17),
    I19   => I(18),
    I20   => I(19),
    I21   => I(20),
    I22   => I(21),
    I23   => I(22),
    I24   => I(23),
    I25   => I(24),
    I26   => I(25),
    I27   => I(26),
    I28   => I(27),
    I29   => I(28),
    I30   => I(29),
    I31   => I(30),
    I32   => I(31),
    I33   => I(32),
    I34   => I(33),
    I35   => I(34),
    I36   => I(35),
    O1    => O(0),
    O2    => O(1),
    O3    => O(2),
    O4    => O(3),
    O5    => O(4),
    O6    => O(5),
    O7    => O(6),
    O8    => O(7),
    O9    => O(8),
    O10   => O(9),
    O11   => O(10),
    O12   => O(11),
    O13   => O(12),
    O14   => O(13),
    O15   => O(14),
    O16   => O(15),
    O17   => O(16),
    O18   => O(17),
    O19   => O(18),
    O20   => O(19),
    O21   => O(20),
    O22   => O(21),
    O23   => O(22),
    O24   => O(23),
    O25   => O(24),
    O26   => O(25),
    O27   => O(26),
    O28   => O(27),
    O29   => O(28),
    O30   => O(29),
    O31   => O(30),
    O32   => O(31),
    O33   => O(32),
    O34   => O(33),
    O35   => O(34),
    O36   => O(35),
    WRSTI => WRSTI,
    WAI1  => WAI(0),
    WAI2  => WAI(1),
    WAI3  => WAI(2),
    WAI4  => WAI(3),
    WAI5  => WAI(4),
    WAI6  => WAI(5),
    WAI7  => '0',
    WAO1  => WAO(0),
    WAO2  => WAO(1),
    WAO3  => WAO(2),
    WAO4  => WAO(3),
    WAO5  => WAO(4),
    WAO6  => WAO(5),
    WAO7  => OPEN,
    WEQ1  => WEQ,
    WEQ2  => OPEN,
    RRSTI => RRSTI,
    RAI1  => RAI(0),
    RAI2  => RAI(1),
    RAI3  => RAI(2),
    RAI4  => RAI(3),
    RAI5  => RAI(4),
    RAI6  => RAI(5),
    RAI7  => '0',
    RAO1  => RAO(0),
    RAO2  => RAO(1),
    RAO3  => RAO(2),
    RAO4  => RAO(3),
    RAO5  => RAO(4),
    RAO6  => RAO(5),
    RAO7  => OPEN,
    REQ1  => REQ,
    REQ2  => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_FIFO_U definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_FIFO_U is
generic (
    mode           : integer := 0; -- 0: DPREG - 1: XFIFO_64x18 - 2: XFIFO_32x36
    wck_edge       : bit := '0';
    rck_edge       : bit := '0';
    use_write_arst : bit := '0';
    use_read_arst  : bit := '0';
    read_addr_inv  : bit_vector(6 downto 0) := "0000000"
);
port (
    RCK    : in  std_logic;
    WCK    : in  std_logic;
    WE     : in  std_logic;
    WEA    : in  std_logic;
    I1     : in  std_logic;
    I2     : in  std_logic;
    I3     : in  std_logic;
    I4     : in  std_logic;
    I5     : in  std_logic;
    I6     : in  std_logic;
    I7     : in  std_logic;
    I8     : in  std_logic;
    I9     : in  std_logic;
    I10    : in  std_logic;
    I11    : in  std_logic;
    I12    : in  std_logic;
    I13    : in  std_logic;
    I14    : in  std_logic;
    I15    : in  std_logic;
    I16    : in  std_logic;
    I17    : in  std_logic;
    I18    : in  std_logic;
    I19    : in  std_logic;
    I20    : in  std_logic;
    I21    : in  std_logic;
    I22    : in  std_logic;
    I23    : in  std_logic;
    I24    : in  std_logic;
    I25    : in  std_logic;
    I26    : in  std_logic;
    I27    : in  std_logic;
    I28    : in  std_logic;
    I29    : in  std_logic;
    I30    : in  std_logic;
    I31    : in  std_logic;
    I32    : in  std_logic;
    I33    : in  std_logic;
    I34    : in  std_logic;
    I35    : in  std_logic;
    I36    : in  std_logic;
    O1     : out std_logic;
    O2     : out std_logic;
    O3     : out std_logic;
    O4     : out std_logic;
    O5     : out std_logic;
    O6     : out std_logic;
    O7     : out std_logic;
    O8     : out std_logic;
    O9     : out std_logic;
    O10    : out std_logic;
    O11    : out std_logic;
    O12    : out std_logic;
    O13    : out std_logic;
    O14    : out std_logic;
    O15    : out std_logic;
    O16    : out std_logic;
    O17    : out std_logic;
    O18    : out std_logic;
    O19    : out std_logic;
    O20    : out std_logic;
    O21    : out std_logic;
    O22    : out std_logic;
    O23    : out std_logic;
    O24    : out std_logic;
    O25    : out std_logic;
    O26    : out std_logic;
    O27    : out std_logic;
    O28    : out std_logic;
    O29    : out std_logic;
    O30    : out std_logic;
    O31    : out std_logic;
    O32    : out std_logic;
    O33    : out std_logic;
    O34    : out std_logic;
    O35    : out std_logic;
    O36    : out std_logic;
    WRSTI  : in  std_logic;
    WAI1   : in  std_logic;
    WAI2   : in  std_logic;
    WAI3   : in  std_logic;
    WAI4   : in  std_logic;
    WAI5   : in  std_logic;
    WAI6   : in  std_logic;
    WAI7   : in  std_logic;
    WAO1   : out std_logic;
    WAO2   : out std_logic;
    WAO3   : out std_logic;
    WAO4   : out std_logic;
    WAO5   : out std_logic;
    WAO6   : out std_logic;
    WAO7   : out std_logic;
    WEQ1   : out std_logic;
    WEQ2   : out std_logic;
    RRSTI  : in  std_logic;
    RAI1   : in  std_logic;
    RAI2   : in  std_logic;
    RAI3   : in  std_logic;
    RAI4   : in  std_logic;
    RAI5   : in  std_logic;
    RAI6   : in  std_logic;
    RAI7   : in  std_logic;
    RAO1   : out std_logic;
    RAO2   : out std_logic;
    RAO3   : out std_logic;
    RAO4   : out std_logic;
    RAO5   : out std_logic;
    RAO6   : out std_logic;
    RAO7   : out std_logic;
    REQ1   : out std_logic;
    REQ2   : out std_logic
);
end NX_FIFO_U;
-- =================================================================================================
--   NX_GCK_U (compatible) definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_GCK_U is
generic (
    inv_in   : bit    := '0';
    inv_out  : bit    := '0';
    std_mode : string := "BYPASS" -- MUX / CKS / BYPASS / CSC
);
port (
    SI1 : in std_logic;
    SI2 : in std_logic;
    CMD : in std_logic;
    SO : out std_logic
);
end NX_GCK_U;
-- =================================================================================================
--   NX_CRX_L definition                                                                2018/11/30
-- =================================================================================================

-- NX_CRX_L#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CRX_L is
 generic (
     test                         : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc           : bit := '0';
     pcs_bypass_usr_cdc           : bit := '0';
     pcs_debug_en                 : bit := '0';
     pcs_fsm_watchdog_en          : bit := '0';
     pma_clk_pos                  : bit := '0';
     pcs_protocol_size            : bit := '0';
     pcs_loopback                 : bit := '0';
     pcs_polarity                 : bit := '0';
     pcs_p_comma_en               : bit := '0';
     pcs_p_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_m_comma_en               : bit := '0';
     pcs_m_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_comma_mask               : bit_vector(9 downto 0) := (others => '0');
     pcs_nb_comma_bef_realign     : bit_vector(1 downto 0) := (others => '0');
     pcs_align_bypass             : bit := '0';
     pcs_dec_bypass               : bit := '0';
     pcs_el_buff_max_comp         : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_diff_bef_comp    : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_only_one_skp     : bit := '0';
     pcs_el_buff_underflow_handle : bit := '0';
     pcs_el_buff_skp_seq_size     : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_char_0       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_1       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_2       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_3       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_size  : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_header_0     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_1     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_2     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_3     : bit_vector(8 downto 0) := (others => '0');
     pcs_buffers_use_cdc          : bit := '0';
     pcs_buffers_bypass           : bit := '0';
     pcs_sync_supported           : bit := '0';
     pcs_replace_bypass           : bit := '0';
     pcs_dscr_bypass              : bit := '0';
     pcs_8b_dscr_sel              : bit := '0';
     pcs_fsm_sel                  : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divf_en_n            : bit := '0';
     pma_pll_divm_en_n            : bit := '0';
     pma_pll_divn_en_n            : bit := '0';
     pma_cdr_cp                   : bit_vector(3 downto 0) := (others => '0');
     pma_ctrl_term                : bit_vector(5 downto 0) := (others => '0');
     pma_pll_cpump_n              : bit_vector(2 downto 0) := (others => '0');
     pma_pll_divf                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divm                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divn                 : bit := '0';
     pma_loopback                 : bit := '0';
     location                     : string := ""
 );
port (
    DSCR_E_I  : in  std_logic;
    DEC_E_I   : in  std_logic;
    ALIGN_E_I : in  std_logic;
    ALIGN_S_I : in  std_logic;
    REP_E_I   : in  std_logic;
    BUF_R_I   : in  std_logic;

    OVS_BS_I1 : in  std_logic;
    OVS_BS_I2 : in  std_logic;

    BUF_FE_I  : in  std_logic;
    RST_N_I   : in  std_logic;
    CDR_R_I   : in  std_logic;
    CKG_RN_I  : in  std_logic;
    PLL_RN_I  : in  std_logic;

    TST_I1    : in  std_logic;
    TST_I2    : in  std_logic;
    TST_I3    : in  std_logic;
    TST_I4    : in  std_logic;

    LOS_O     : out std_logic;

    DATA_O1   : out std_logic;
    DATA_O2   : out std_logic;
    DATA_O3   : out std_logic;
    DATA_O4   : out std_logic;
    DATA_O5   : out std_logic;
    DATA_O6   : out std_logic;
    DATA_O7   : out std_logic;
    DATA_O8   : out std_logic;
    DATA_O9   : out std_logic;
    DATA_O10  : out std_logic;
    DATA_O11  : out std_logic;
    DATA_O12  : out std_logic;
    DATA_O13  : out std_logic;
    DATA_O14  : out std_logic;
    DATA_O15  : out std_logic;
    DATA_O16  : out std_logic;
    DATA_O17  : out std_logic;
    DATA_O18  : out std_logic;
    DATA_O19  : out std_logic;
    DATA_O20  : out std_logic;
    DATA_O21  : out std_logic;
    DATA_O22  : out std_logic;
    DATA_O23  : out std_logic;
    DATA_O24  : out std_logic;
    DATA_O25  : out std_logic;
    DATA_O26  : out std_logic;
    DATA_O27  : out std_logic;
    DATA_O28  : out std_logic;
    DATA_O29  : out std_logic;
    DATA_O30  : out std_logic;
    DATA_O31  : out std_logic;
    DATA_O32  : out std_logic;
    DATA_O33  : out std_logic;
    DATA_O34  : out std_logic;
    DATA_O35  : out std_logic;
    DATA_O36  : out std_logic;
    DATA_O37  : out std_logic;
    DATA_O38  : out std_logic;
    DATA_O39  : out std_logic;
    DATA_O40  : out std_logic;
    DATA_O41  : out std_logic;
    DATA_O42  : out std_logic;
    DATA_O43  : out std_logic;
    DATA_O44  : out std_logic;
    DATA_O45  : out std_logic;
    DATA_O46  : out std_logic;
    DATA_O47  : out std_logic;
    DATA_O48  : out std_logic;
    DATA_O49  : out std_logic;
    DATA_O50  : out std_logic;
    DATA_O51  : out std_logic;
    DATA_O52  : out std_logic;
    DATA_O53  : out std_logic;
    DATA_O54  : out std_logic;
    DATA_O55  : out std_logic;
    DATA_O56  : out std_logic;
    DATA_O57  : out std_logic;
    DATA_O58  : out std_logic;
    DATA_O59  : out std_logic;
    DATA_O60  : out std_logic;
    DATA_O61  : out std_logic;
    DATA_O62  : out std_logic;
    DATA_O63  : out std_logic;
    DATA_O64  : out std_logic;

    CH_COM_O1 : out std_logic;
    CH_COM_O2 : out std_logic;
    CH_COM_O3 : out std_logic;
    CH_COM_O4 : out std_logic;
    CH_COM_O5 : out std_logic;
    CH_COM_O6 : out std_logic;
    CH_COM_O7 : out std_logic;
    CH_COM_O8 : out std_logic;

    CH_K_O1   : out std_logic;
    CH_K_O2   : out std_logic;
    CH_K_O3   : out std_logic;
    CH_K_O4   : out std_logic;
    CH_K_O5   : out std_logic;
    CH_K_O6   : out std_logic;
    CH_K_O7   : out std_logic;
    CH_K_O8   : out std_logic;

    NIT_O1    : out std_logic;
    NIT_O2    : out std_logic;
    NIT_O3    : out std_logic;
    NIT_O4    : out std_logic;
    NIT_O5    : out std_logic;
    NIT_O6    : out std_logic;
    NIT_O7    : out std_logic;
    NIT_O8    : out std_logic;

    D_ERR_O1  : out std_logic;
    D_ERR_O2  : out std_logic;
    D_ERR_O3  : out std_logic;
    D_ERR_O4  : out std_logic;
    D_ERR_O5  : out std_logic;
    D_ERR_O6  : out std_logic;
    D_ERR_O7  : out std_logic;
    D_ERR_O8  : out std_logic;

    CH_A_O1   : out std_logic;
    CH_A_O2   : out std_logic;
    CH_A_O3   : out std_logic;
    CH_A_O4   : out std_logic;
    CH_A_O5   : out std_logic;
    CH_A_O6   : out std_logic;
    CH_A_O7   : out std_logic;
    CH_A_O8   : out std_logic;

    CH_F_O1   : out std_logic;
    CH_F_O2   : out std_logic;
    CH_F_O3   : out std_logic;
    CH_F_O4   : out std_logic;
    CH_F_O5   : out std_logic;
    CH_F_O6   : out std_logic;
    CH_F_O7   : out std_logic;
    CH_F_O8   : out std_logic;

    ALIGN_O   : out std_logic;
    BUSY_O    : out std_logic;

    TST_O1    : out std_logic;
    TST_O2    : out std_logic;
    TST_O3    : out std_logic;
    TST_O4    : out std_logic;
    TST_O5    : out std_logic;
    TST_O6    : out std_logic;
    TST_O7    : out std_logic;
    TST_O8    : out std_logic;

    LOCK_O    : out std_logic;

    LINK      : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);

    RX_I      : in  std_logic
);
end NX_CRX_L;
--#}}}#
-- =================================================================================================
--   NX_CTX_L definition                                                                2018/11/30
-- =================================================================================================

-- NX_CTX_L#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CTX_L is
 generic (
     pma_clk_pos          : bit := '0';
     pcs_protocol_size    : bit := '0';
     pcs_8b_scr_sel       : bit := '0';
     pcs_scr_init         : bit_vector(16 downto 0) := (others => '0');
     pcs_scr_bypass       : bit := '0';
     pcs_sync_supported   : bit := '0';
     pcs_replace_bypass   : bit := '0';
     pcs_enc_bypass       : bit := '0';
     pcs_loopback         : bit := '0';
     pcs_polarity         : bit := '0';
     pcs_esistream_fsm_en : bit := '0';
     test                 : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc   : bit := '0';
     pcs_bypass_usr_cdc   : bit := '0';
     pma_loopback         : bit := '0';
     location             : string := ""
 );
port (
    ENC_E_I1 : in  std_logic;
    ENC_E_I2 : in  std_logic;
    ENC_E_I3 : in  std_logic;
    ENC_E_I4 : in  std_logic;
    ENC_E_I5 : in  std_logic;
    ENC_E_I6 : in  std_logic;
    ENC_E_I7 : in  std_logic;
    ENC_E_I8 : in  std_logic;

    CH_K_I1  : in  std_logic;
    CH_K_I2  : in  std_logic;
    CH_K_I3  : in  std_logic;
    CH_K_I4  : in  std_logic;
    CH_K_I5  : in  std_logic;
    CH_K_I6  : in  std_logic;
    CH_K_I7  : in  std_logic;
    CH_K_I8  : in  std_logic;

    SCR_E_I1 : in  std_logic;
    SCR_E_I2 : in  std_logic;
    SCR_E_I3 : in  std_logic;
    SCR_E_I4 : in  std_logic;
    SCR_E_I5 : in  std_logic;
    SCR_E_I6 : in  std_logic;
    SCR_E_I7 : in  std_logic;
    SCR_E_I8 : in  std_logic;

    EOMF_I1  : in  std_logic;
    EOMF_I2  : in  std_logic;
    EOMF_I3  : in  std_logic;
    EOMF_I4  : in  std_logic;
    EOMF_I5  : in  std_logic;
    EOMF_I6  : in  std_logic;
    EOMF_I7  : in  std_logic;
    EOMF_I8  : in  std_logic;

    EOF_I1   : in  std_logic;
    EOF_I2   : in  std_logic;
    EOF_I3   : in  std_logic;
    EOF_I4   : in  std_logic;
    EOF_I5   : in  std_logic;
    EOF_I6   : in  std_logic;
    EOF_I7   : in  std_logic;
    EOF_I8   : in  std_logic;

    REP_E_I  : in  std_logic;
    RST_N_I  : in  std_logic;

    TST_I1   : in  std_logic;
    TST_I2   : in  std_logic;
    TST_I3   : in  std_logic;
    TST_I4   : in  std_logic;

    DATA_I1  : in  std_logic;
    DATA_I2  : in  std_logic;
    DATA_I3  : in  std_logic;
    DATA_I4  : in  std_logic;
    DATA_I5  : in  std_logic;
    DATA_I6  : in  std_logic;
    DATA_I7  : in  std_logic;
    DATA_I8  : in  std_logic;
    DATA_I9  : in  std_logic;
    DATA_I10 : in  std_logic;
    DATA_I11 : in  std_logic;
    DATA_I12 : in  std_logic;
    DATA_I13 : in  std_logic;
    DATA_I14 : in  std_logic;
    DATA_I15 : in  std_logic;
    DATA_I16 : in  std_logic;
    DATA_I17 : in  std_logic;
    DATA_I18 : in  std_logic;
    DATA_I19 : in  std_logic;
    DATA_I20 : in  std_logic;
    DATA_I21 : in  std_logic;
    DATA_I22 : in  std_logic;
    DATA_I23 : in  std_logic;
    DATA_I24 : in  std_logic;
    DATA_I25 : in  std_logic;
    DATA_I26 : in  std_logic;
    DATA_I27 : in  std_logic;
    DATA_I28 : in  std_logic;
    DATA_I29 : in  std_logic;
    DATA_I30 : in  std_logic;
    DATA_I31 : in  std_logic;
    DATA_I32 : in  std_logic;
    DATA_I33 : in  std_logic;
    DATA_I34 : in  std_logic;
    DATA_I35 : in  std_logic;
    DATA_I36 : in  std_logic;
    DATA_I37 : in  std_logic;
    DATA_I38 : in  std_logic;
    DATA_I39 : in  std_logic;
    DATA_I40 : in  std_logic;
    DATA_I41 : in  std_logic;
    DATA_I42 : in  std_logic;
    DATA_I43 : in  std_logic;
    DATA_I44 : in  std_logic;
    DATA_I45 : in  std_logic;
    DATA_I46 : in  std_logic;
    DATA_I47 : in  std_logic;
    DATA_I48 : in  std_logic;
    DATA_I49 : in  std_logic;
    DATA_I50 : in  std_logic;
    DATA_I51 : in  std_logic;
    DATA_I52 : in  std_logic;
    DATA_I53 : in  std_logic;
    DATA_I54 : in  std_logic;
    DATA_I55 : in  std_logic;
    DATA_I56 : in  std_logic;
    DATA_I57 : in  std_logic;
    DATA_I58 : in  std_logic;
    DATA_I59 : in  std_logic;
    DATA_I60 : in  std_logic;
    DATA_I61 : in  std_logic;
    DATA_I62 : in  std_logic;
    DATA_I63 : in  std_logic;
    DATA_I64 : in  std_logic;

    TST_O1   : out std_logic;
    TST_O2   : out std_logic;
    TST_O3   : out std_logic;
    TST_O4   : out std_logic;

    BUSY_O   : out std_logic;
    CLK_E_I  : in  std_logic;

    LINK     : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);

    TX_O     : out std_logic
);
end NX_CTX_L;
--#}}}#
-- =================================================================================================
--   NX_HSSL_L_FULL declaration                                                          2019/06/20
-- =================================================================================================

-- NX_HSSL_L_FULL#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_HSSL_L_FULL is
generic (
   cfg_main_i : bit_vector( 33 downto 0) := (others => '0');
   cfg_tx0_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx0_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx1_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx1_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx2_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx2_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx3_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx3_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx4_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx4_i  : bit_vector(159 downto 0) := (others => '0');
   cfg_tx5_i  : bit_vector( 31 downto 0) := (others => '0');
   cfg_rx5_i  : bit_vector(159 downto 0) := (others => '0');
   location   : string := ""
 );
port (
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ MAIN ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- Fabric Interface
   hssl_clk_user_i                       : in  std_logic;
   hssl_clk_ref_i                        : in  std_logic;
   hssl_clock_o                          : out std_logic;
   usr_com_tx_pma_pre_sign_i             : in  std_logic;
   usr_com_tx_pma_pre_en_i               : in  std_logic;
   usr_com_tx_pma_pre_input_sel_i        : in  std_logic_vector(3 downto 0);
   usr_com_tx_pma_main_sign_i            : in  std_logic;
   usr_com_rx_pma_m_eye_i                : in  std_logic;
   usr_com_tx_pma_main_en_i              : in  std_logic_vector(5 downto 0);
   usr_com_tx_pma_margin_sel_i           : in  std_logic_vector(3 downto 0);
   usr_com_tx_pma_margin_input_sel_i     : in  std_logic_vector(3 downto 0);
   usr_com_tx_pma_margin_sel_var_i       : in  std_logic_vector(4 downto 0);
   usr_com_tx_pma_margin_input_sel_var_i : in  std_logic_vector(4 downto 0);
   usr_com_tx_pma_post_en_i              : in  std_logic_vector(4 downto 0);
   usr_com_tx_pma_post_sign_i            : in  std_logic;
   usr_com_tx_pma_post_input_sel_i       : in  std_logic_vector(3 downto 0);
   usr_com_tx_pma_post_input_sel_var_i   : in  std_logic_vector(3 downto 0);
   usr_com_rx_pma_ctle_cap_i             : in  std_logic_vector(3 downto 0);
   usr_com_rx_pma_ctle_resp_i            : in  std_logic_vector(3 downto 0);
   usr_com_rx_pma_ctle_resn_i            : in  std_logic_vector(3 downto 0);
   usr_com_ctrl_tx_sel_i                 : in  std_logic_vector(5 downto 0);
   usr_com_ctrl_rx_sel_i                 : in  std_logic_vector(5 downto 0);
   usr_pll_pma_rst_n_i                   : in  std_logic;
   usr_main_rst_n_i                      : in  std_logic;
   usr_calibrate_pma_res_p1_i            : in  std_logic_vector(7 downto 0);
   usr_calibrate_pma_res_n2_i            : in  std_logic_vector(7 downto 0);
   usr_calibrate_pma_res_n3_i            : in  std_logic_vector(7 downto 0);
   usr_calibrate_pma_res_p4_i            : in  std_logic_vector(7 downto 0);
   usr_calibrate_pma_sel_i               : in  std_logic_vector(3 downto 0);
   usr_calibrate_pma_en_i                : in  std_logic;
   usr_pcs_ctrl_pll_lock_en_i            : in  std_logic;
   usr_pcs_ctrl_ovs_en_i                 : in  std_logic;
   usr_main_test_i                       : in  std_logic_vector(7 downto 0);
   usr_pll_lock_o                        : out std_logic;
   usr_calibrate_pma_out_o               : out std_logic;
   usr_main_test_o                       : out std_logic_vector(7 downto 0);
   pma_clk_ext_i                         : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 0 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx0_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_replace_en_i        : in  std_logic;
   usr_tx0_rst_n_i                  : in  std_logic;
   usr_tx0_pma_clk_en_i             : in  std_logic;
   usr_tx0_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx0_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx0_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx0_busy_o                   : out std_logic;
   pma_tx0_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx0_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx0_ctrl_dscr_en_i         : in  std_logic;
   usr_rx0_ctrl_dec_en_i          : in  std_logic;
   usr_rx0_ctrl_align_en_i        : in  std_logic;
   usr_rx0_ctrl_align_sync_i      : in  std_logic;
   usr_rx0_ctrl_replace_en_i      : in  std_logic;
   usr_rx0_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx0_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx0_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx0_rst_n_i                : in  std_logic;
   usr_rx0_pma_cdr_rst_i          : in  std_logic;
   usr_rx0_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx0_pma_pll_rst_n_i        : in  std_logic;
   usr_rx0_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx0_pma_loss_of_signal_o   : out std_logic;
   usr_rx0_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_aligned_o : out std_logic;
   usr_rx0_busy_o                 : out std_logic;
   usr_rx0_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx0_pll_lock_o             : out std_logic;
   pma_rx0_i                      : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 1 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx1_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_replace_en_i        : in  std_logic;
   usr_tx1_rst_n_i                  : in  std_logic;
   usr_tx1_pma_clk_en_i             : in  std_logic;
   usr_tx1_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx1_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx1_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx1_busy_o                   : out std_logic;
   pma_tx1_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx1_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx1_ctrl_dscr_en_i         : in  std_logic;
   usr_rx1_ctrl_dec_en_i          : in  std_logic;
   usr_rx1_ctrl_align_en_i        : in  std_logic;
   usr_rx1_ctrl_align_sync_i      : in  std_logic;
   usr_rx1_ctrl_replace_en_i      : in  std_logic;
   usr_rx1_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx1_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx1_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx1_rst_n_i                : in  std_logic;
   usr_rx1_pma_cdr_rst_i          : in  std_logic;
   usr_rx1_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx1_pma_pll_rst_n_i        : in  std_logic;
   usr_rx1_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx1_pma_loss_of_signal_o   : out std_logic;
   usr_rx1_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_aligned_o : out std_logic;
   usr_rx1_busy_o                 : out std_logic;
   usr_rx1_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx1_pll_lock_o             : out std_logic;
   pma_rx1_i                      : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 2 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx2_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_replace_en_i        : in  std_logic;
   usr_tx2_rst_n_i                  : in  std_logic;
   usr_tx2_pma_clk_en_i             : in  std_logic;
   usr_tx2_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx2_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx2_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx2_busy_o                   : out std_logic;
   pma_tx2_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx2_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx2_ctrl_dscr_en_i         : in  std_logic;
   usr_rx2_ctrl_dec_en_i          : in  std_logic;
   usr_rx2_ctrl_align_en_i        : in  std_logic;
   usr_rx2_ctrl_align_sync_i      : in  std_logic;
   usr_rx2_ctrl_replace_en_i      : in  std_logic;
   usr_rx2_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx2_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx2_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx2_rst_n_i                : in  std_logic;
   usr_rx2_pma_cdr_rst_i          : in  std_logic;
   usr_rx2_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx2_pma_pll_rst_n_i        : in  std_logic;
   usr_rx2_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx2_pma_loss_of_signal_o   : out std_logic;
   usr_rx2_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_aligned_o : out std_logic;
   usr_rx2_busy_o                 : out std_logic;
   usr_rx2_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx2_pll_lock_o             : out std_logic;
   pma_rx2_i                      : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 3 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx3_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_replace_en_i        : in  std_logic;
   usr_tx3_rst_n_i                  : in  std_logic;
   usr_tx3_pma_clk_en_i             : in  std_logic;
   usr_tx3_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx3_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx3_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx3_busy_o                   : out std_logic;
   pma_tx3_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx3_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx3_ctrl_dscr_en_i         : in  std_logic;
   usr_rx3_ctrl_dec_en_i          : in  std_logic;
   usr_rx3_ctrl_align_en_i        : in  std_logic;
   usr_rx3_ctrl_align_sync_i      : in  std_logic;
   usr_rx3_ctrl_replace_en_i      : in  std_logic;
   usr_rx3_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx3_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx3_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx3_rst_n_i                : in  std_logic;
   usr_rx3_pma_cdr_rst_i          : in  std_logic;
   usr_rx3_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx3_pma_pll_rst_n_i        : in  std_logic;
   usr_rx3_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx3_pma_loss_of_signal_o   : out std_logic;
   usr_rx3_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_aligned_o : out std_logic;
   usr_rx3_busy_o                 : out std_logic;
   usr_rx3_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx3_pll_lock_o             : out std_logic;
   pma_rx3_i                      : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 4 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx4_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx4_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx4_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx4_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx4_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx4_ctrl_replace_en_i        : in  std_logic;
   usr_tx4_rst_n_i                  : in  std_logic;
   usr_tx4_pma_clk_en_i             : in  std_logic;
   usr_tx4_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx4_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx4_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx4_busy_o                   : out std_logic;
   pma_tx4_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx4_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx4_ctrl_dscr_en_i         : in  std_logic;
   usr_rx4_ctrl_dec_en_i          : in  std_logic;
   usr_rx4_ctrl_align_en_i        : in  std_logic;
   usr_rx4_ctrl_align_sync_i      : in  std_logic;
   usr_rx4_ctrl_replace_en_i      : in  std_logic;
   usr_rx4_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx4_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx4_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx4_rst_n_i                : in  std_logic;
   usr_rx4_pma_cdr_rst_i          : in  std_logic;
   usr_rx4_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx4_pma_pll_rst_n_i        : in  std_logic;
   usr_rx4_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx4_pma_loss_of_signal_o   : out std_logic;
   usr_rx4_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx4_ctrl_char_is_aligned_o : out std_logic;
   usr_rx4_busy_o                 : out std_logic;
   usr_rx4_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx4_pll_lock_o             : out std_logic;
   pma_rx4_i                      : in  std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 5 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
    -- TX - Fabric Interface
   usr_tx5_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx5_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx5_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx5_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx5_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx5_ctrl_replace_en_i        : in  std_logic;
   usr_tx5_rst_n_i                  : in  std_logic;
   usr_tx5_pma_clk_en_i             : in  std_logic;
   usr_tx5_test_i                   : in  std_logic_vector(3 downto 0);
   usr_tx5_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx5_test_o                   : out std_logic_vector(3 downto 0);
   usr_tx5_busy_o                   : out std_logic;
   pma_tx5_o                        : out std_logic;
    -- RX - Fabric Interface
   usr_rx5_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx5_ctrl_dscr_en_i         : in  std_logic;
   usr_rx5_ctrl_dec_en_i          : in  std_logic;
   usr_rx5_ctrl_align_en_i        : in  std_logic;
   usr_rx5_ctrl_align_sync_i      : in  std_logic;
   usr_rx5_ctrl_replace_en_i      : in  std_logic;
   usr_rx5_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx5_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx5_ctrl_el_buff_fifo_en_i : in  std_logic;
   usr_rx5_rst_n_i                : in  std_logic;
   usr_rx5_pma_cdr_rst_i          : in  std_logic;
   usr_rx5_pma_ckgen_rst_n_i      : in  std_logic;
   usr_rx5_pma_pll_rst_n_i        : in  std_logic;
   usr_rx5_test_i                 : in  std_logic_vector(3 downto 0);
   usr_rx5_pma_loss_of_signal_o   : out std_logic;
   usr_rx5_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx5_ctrl_char_is_aligned_o : out std_logic;
   usr_rx5_busy_o                 : out std_logic;
   usr_rx5_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx5_pll_lock_o             : out std_logic;
   pma_rx5_i                      : in  std_logic
);
end NX_HSSL_L_FULL;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_HSSL_L_FULL definition                                                           2019/06/20
-- =================================================================================================

-- NX_HSSL_L_FULL#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

architecture NX_RTL of NX_HSSL_L_FULL is

signal LINK_RX0 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX1 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX2 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX3 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX4 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX5 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_TX0 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX1 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX2 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX3 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX4 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX5 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);

-- component NX_CTX_L#{{{#
component NX_CTX_L
 generic (
     pma_clk_pos          : bit := '0';
     pcs_protocol_size    : bit := '0';
     pcs_8b_scr_sel       : bit := '0';
     pcs_scr_init         : bit_vector(16 downto 0) := (others => '0');
     pcs_scr_bypass       : bit := '0';
     pcs_sync_supported   : bit := '0';
     pcs_replace_bypass   : bit := '0';
     pcs_loopback         : bit := '0';
     pcs_enc_bypass       : bit := '0';
     pcs_polarity         : bit := '0';
     pcs_esistream_fsm_en : bit := '0';
     test                 : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc   : bit := '0';
     pcs_bypass_usr_cdc   : bit := '0';
     pma_loopback         : bit := '0';
     location             : string := ""
 );
port (
    ENC_E_I1 : in  std_logic;
    ENC_E_I2 : in  std_logic;
    ENC_E_I3 : in  std_logic;
    ENC_E_I4 : in  std_logic;
    ENC_E_I5 : in  std_logic;
    ENC_E_I6 : in  std_logic;
    ENC_E_I7 : in  std_logic;
    ENC_E_I8 : in  std_logic;

    CH_K_I1  : in  std_logic;
    CH_K_I2  : in  std_logic;
    CH_K_I3  : in  std_logic;
    CH_K_I4  : in  std_logic;
    CH_K_I5  : in  std_logic;
    CH_K_I6  : in  std_logic;
    CH_K_I7  : in  std_logic;
    CH_K_I8  : in  std_logic;

    SCR_E_I1 : in  std_logic;
    SCR_E_I2 : in  std_logic;
    SCR_E_I3 : in  std_logic;
    SCR_E_I4 : in  std_logic;
    SCR_E_I5 : in  std_logic;
    SCR_E_I6 : in  std_logic;
    SCR_E_I7 : in  std_logic;
    SCR_E_I8 : in  std_logic;

    EOMF_I1  : in  std_logic;
    EOMF_I2  : in  std_logic;
    EOMF_I3  : in  std_logic;
    EOMF_I4  : in  std_logic;
    EOMF_I5  : in  std_logic;
    EOMF_I6  : in  std_logic;
    EOMF_I7  : in  std_logic;
    EOMF_I8  : in  std_logic;

    EOF_I1   : in  std_logic;
    EOF_I2   : in  std_logic;
    EOF_I3   : in  std_logic;
    EOF_I4   : in  std_logic;
    EOF_I5   : in  std_logic;
    EOF_I6   : in  std_logic;
    EOF_I7   : in  std_logic;
    EOF_I8   : in  std_logic;

    REP_E_I  : in  std_logic;
    RST_N_I  : in  std_logic;

    TST_I1   : in  std_logic;
    TST_I2   : in  std_logic;
    TST_I3   : in  std_logic;
    TST_I4   : in  std_logic;

    DATA_I1  : in  std_logic;
    DATA_I2  : in  std_logic;
    DATA_I3  : in  std_logic;
    DATA_I4  : in  std_logic;
    DATA_I5  : in  std_logic;
    DATA_I6  : in  std_logic;
    DATA_I7  : in  std_logic;
    DATA_I8  : in  std_logic;
    DATA_I9  : in  std_logic;
    DATA_I10 : in  std_logic;
    DATA_I11 : in  std_logic;
    DATA_I12 : in  std_logic;
    DATA_I13 : in  std_logic;
    DATA_I14 : in  std_logic;
    DATA_I15 : in  std_logic;
    DATA_I16 : in  std_logic;
    DATA_I17 : in  std_logic;
    DATA_I18 : in  std_logic;
    DATA_I19 : in  std_logic;
    DATA_I20 : in  std_logic;
    DATA_I21 : in  std_logic;
    DATA_I22 : in  std_logic;
    DATA_I23 : in  std_logic;
    DATA_I24 : in  std_logic;
    DATA_I25 : in  std_logic;
    DATA_I26 : in  std_logic;
    DATA_I27 : in  std_logic;
    DATA_I28 : in  std_logic;
    DATA_I29 : in  std_logic;
    DATA_I30 : in  std_logic;
    DATA_I31 : in  std_logic;
    DATA_I32 : in  std_logic;
    DATA_I33 : in  std_logic;
    DATA_I34 : in  std_logic;
    DATA_I35 : in  std_logic;
    DATA_I36 : in  std_logic;
    DATA_I37 : in  std_logic;
    DATA_I38 : in  std_logic;
    DATA_I39 : in  std_logic;
    DATA_I40 : in  std_logic;
    DATA_I41 : in  std_logic;
    DATA_I42 : in  std_logic;
    DATA_I43 : in  std_logic;
    DATA_I44 : in  std_logic;
    DATA_I45 : in  std_logic;
    DATA_I46 : in  std_logic;
    DATA_I47 : in  std_logic;
    DATA_I48 : in  std_logic;
    DATA_I49 : in  std_logic;
    DATA_I50 : in  std_logic;
    DATA_I51 : in  std_logic;
    DATA_I52 : in  std_logic;
    DATA_I53 : in  std_logic;
    DATA_I54 : in  std_logic;
    DATA_I55 : in  std_logic;
    DATA_I56 : in  std_logic;
    DATA_I57 : in  std_logic;
    DATA_I58 : in  std_logic;
    DATA_I59 : in  std_logic;
    DATA_I60 : in  std_logic;
    DATA_I61 : in  std_logic;
    DATA_I62 : in  std_logic;
    DATA_I63 : in  std_logic;
    DATA_I64 : in  std_logic;

    TST_O1   : out std_logic;
    TST_O2   : out std_logic;
    TST_O3   : out std_logic;
    TST_O4   : out std_logic;

    BUSY_O   : out std_logic;
    CLK_E_I  : in  std_logic;

    LINK     : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);

    TX_O     : out std_logic
);
end component;
--#}}}#

-- component NX_CRX_L#{{{#
component NX_CRX_L
 generic (
     test                         : bit_vector(1 downto 0) := (others => '0');
     pcs_bypass_pma_cdc           : bit := '0';
     pcs_bypass_usr_cdc           : bit := '0';
     pcs_debug_en                 : bit := '0';
     pcs_fsm_watchdog_en          : bit := '0';
     pma_clk_pos                  : bit := '0';
     pcs_protocol_size            : bit := '0';
     pcs_loopback                 : bit := '0';
     pcs_polarity                 : bit := '0';
     pcs_p_comma_en               : bit := '0';
     pcs_p_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_m_comma_en               : bit := '0';
     pcs_m_comma_val              : bit_vector(9 downto 0) := (others => '0');
     pcs_comma_mask               : bit_vector(9 downto 0) := (others => '0');
     pcs_nb_comma_bef_realign     : bit_vector(1 downto 0) := (others => '0');
     pcs_align_bypass             : bit := '0';
     pcs_dec_bypass               : bit := '0';
     pcs_el_buff_max_comp         : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_diff_bef_comp    : bit_vector(2 downto 0) := (others => '0');
     pcs_el_buff_only_one_skp     : bit := '0';
     pcs_el_buff_underflow_handle : bit := '0';
     pcs_el_buff_skp_seq_size     : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_char_0       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_1       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_2       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_char_3       : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_size  : bit_vector(1 downto 0) := (others => '0');
     pcs_el_buff_skp_header_0     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_1     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_2     : bit_vector(8 downto 0) := (others => '0');
     pcs_el_buff_skp_header_3     : bit_vector(8 downto 0) := (others => '0');
     pcs_buffers_use_cdc          : bit := '0';
     pcs_buffers_bypass           : bit := '0';
     pcs_sync_supported           : bit := '0';
     pcs_replace_bypass           : bit := '0';
     pcs_dscr_bypass              : bit := '0';
     pcs_8b_dscr_sel              : bit := '0';
     pcs_fsm_sel                  : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divf_en_n            : bit := '0';
     pma_pll_divm_en_n            : bit := '0';
     pma_pll_divn_en_n            : bit := '0';
     pma_cdr_cp                   : bit_vector(3 downto 0) := (others => '0');
     pma_ctrl_term                : bit_vector(5 downto 0) := (others => '0');
     pma_pll_cpump_n              : bit_vector(2 downto 0) := (others => '0');
     pma_pll_divf                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divm                 : bit_vector(1 downto 0) := (others => '0');
     pma_pll_divn                 : bit := '0';
     pma_loopback                 : bit := '0';
     location                     : string := ""
 );
port (
    DSCR_E_I  : in  std_logic;
    DEC_E_I   : in  std_logic;
    ALIGN_E_I : in  std_logic;
    ALIGN_S_I : in  std_logic;
    REP_E_I   : in  std_logic;
    BUF_R_I   : in  std_logic;

    OVS_BS_I1 : in  std_logic;
    OVS_BS_I2 : in  std_logic;

    BUF_FE_I  : in  std_logic;
    RST_N_I   : in  std_logic;
    CDR_R_I   : in  std_logic;
    CKG_RN_I  : in  std_logic;
    PLL_RN_I  : in  std_logic;

    TST_I1    : in  std_logic;
    TST_I2    : in  std_logic;
    TST_I3    : in  std_logic;
    TST_I4    : in  std_logic;

    LOS_O     : out std_logic;

    DATA_O1   : out std_logic;
    DATA_O2   : out std_logic;
    DATA_O3   : out std_logic;
    DATA_O4   : out std_logic;
    DATA_O5   : out std_logic;
    DATA_O6   : out std_logic;
    DATA_O7   : out std_logic;
    DATA_O8   : out std_logic;
    DATA_O9   : out std_logic;
    DATA_O10  : out std_logic;
    DATA_O11  : out std_logic;
    DATA_O12  : out std_logic;
    DATA_O13  : out std_logic;
    DATA_O14  : out std_logic;
    DATA_O15  : out std_logic;
    DATA_O16  : out std_logic;
    DATA_O17  : out std_logic;
    DATA_O18  : out std_logic;
    DATA_O19  : out std_logic;
    DATA_O20  : out std_logic;
    DATA_O21  : out std_logic;
    DATA_O22  : out std_logic;
    DATA_O23  : out std_logic;
    DATA_O24  : out std_logic;
    DATA_O25  : out std_logic;
    DATA_O26  : out std_logic;
    DATA_O27  : out std_logic;
    DATA_O28  : out std_logic;
    DATA_O29  : out std_logic;
    DATA_O30  : out std_logic;
    DATA_O31  : out std_logic;
    DATA_O32  : out std_logic;
    DATA_O33  : out std_logic;
    DATA_O34  : out std_logic;
    DATA_O35  : out std_logic;
    DATA_O36  : out std_logic;
    DATA_O37  : out std_logic;
    DATA_O38  : out std_logic;
    DATA_O39  : out std_logic;
    DATA_O40  : out std_logic;
    DATA_O41  : out std_logic;
    DATA_O42  : out std_logic;
    DATA_O43  : out std_logic;
    DATA_O44  : out std_logic;
    DATA_O45  : out std_logic;
    DATA_O46  : out std_logic;
    DATA_O47  : out std_logic;
    DATA_O48  : out std_logic;
    DATA_O49  : out std_logic;
    DATA_O50  : out std_logic;
    DATA_O51  : out std_logic;
    DATA_O52  : out std_logic;
    DATA_O53  : out std_logic;
    DATA_O54  : out std_logic;
    DATA_O55  : out std_logic;
    DATA_O56  : out std_logic;
    DATA_O57  : out std_logic;
    DATA_O58  : out std_logic;
    DATA_O59  : out std_logic;
    DATA_O60  : out std_logic;
    DATA_O61  : out std_logic;
    DATA_O62  : out std_logic;
    DATA_O63  : out std_logic;
    DATA_O64  : out std_logic;

    CH_COM_O1 : out std_logic;
    CH_COM_O2 : out std_logic;
    CH_COM_O3 : out std_logic;
    CH_COM_O4 : out std_logic;
    CH_COM_O5 : out std_logic;
    CH_COM_O6 : out std_logic;
    CH_COM_O7 : out std_logic;
    CH_COM_O8 : out std_logic;

    CH_K_O1   : out std_logic;
    CH_K_O2   : out std_logic;
    CH_K_O3   : out std_logic;
    CH_K_O4   : out std_logic;
    CH_K_O5   : out std_logic;
    CH_K_O6   : out std_logic;
    CH_K_O7   : out std_logic;
    CH_K_O8   : out std_logic;

    NIT_O1    : out std_logic;
    NIT_O2    : out std_logic;
    NIT_O3    : out std_logic;
    NIT_O4    : out std_logic;
    NIT_O5    : out std_logic;
    NIT_O6    : out std_logic;
    NIT_O7    : out std_logic;
    NIT_O8    : out std_logic;

    D_ERR_O1  : out std_logic;
    D_ERR_O2  : out std_logic;
    D_ERR_O3  : out std_logic;
    D_ERR_O4  : out std_logic;
    D_ERR_O5  : out std_logic;
    D_ERR_O6  : out std_logic;
    D_ERR_O7  : out std_logic;
    D_ERR_O8  : out std_logic;

    CH_A_O1   : out std_logic;
    CH_A_O2   : out std_logic;
    CH_A_O3   : out std_logic;
    CH_A_O4   : out std_logic;
    CH_A_O5   : out std_logic;
    CH_A_O6   : out std_logic;
    CH_A_O7   : out std_logic;
    CH_A_O8   : out std_logic;
    CH_F_O1   : out std_logic;
    CH_F_O2   : out std_logic;
    CH_F_O3   : out std_logic;
    CH_F_O4   : out std_logic;
    CH_F_O5   : out std_logic;
    CH_F_O6   : out std_logic;
    CH_F_O7   : out std_logic;
    CH_F_O8   : out std_logic;

    ALIGN_O   : out std_logic;
    BUSY_O    : out std_logic;

    TST_O1    : out std_logic;
    TST_O2    : out std_logic;
    TST_O3    : out std_logic;
    TST_O4    : out std_logic;
    TST_O5    : out std_logic;
    TST_O6    : out std_logic;
    TST_O7    : out std_logic;
    TST_O8    : out std_logic;

    LOCK_O    : out std_logic;

    LINK      : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);

    RX_I      : in  std_logic
);
end component;
--#}}}#

-- component NX_PMA_L#{{{#
component NX_PMA_L
 generic (
     main_test                   : bit_vector(7 downto 0) := (others => '0');
     rx_pma_half_step            : bit := '0';
     pll_pma_int_data_len        : bit := '0';
     pll_pma_cpump_n             : bit_vector(2 downto 0) := (others => '0');
     pll_pma_divf                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divm                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divn                : bit := '0';
     pll_pma_lvds_mux            : bit := '0';
     pll_pma_mux_ckref           : bit := '0';
     pll_pma_divf_en_n           : bit := '0';
     pll_pma_divm_en_n           : bit := '0';
     pll_pma_divn_en_n           : bit := '0';
     main_clk_to_fabric_div_mode : bit := '0';
     main_clk_to_fabric_div_en   : bit := '0';
     main_clk_to_fabric_sel      : bit := '0';
     main_use_only_usr_clock     : bit := '0';
     main_use_pcs_clk_2          : bit := '0';
     pcs_word_len                : bit_vector(1 downto 0) := (others => '0');
     pcs_ovs_mode                : bit := '0';
     pcs_pll_lock_count          : bit_vector(2 downto 0) := (others => '0');
     location                    : string := ""
 );
port (
    CLK_USER_I  : in  std_logic;
    CLK_REF_I   : in  std_logic;
--    CLK_I1      : in  std_logic;
--    CLK_I2      : in  std_logic;
--    CLK_I3      : in  std_logic;
--    CLK_I4      : in  std_logic;
--    CLK_I5      : in  std_logic;
--    CLK_I6      : in  std_logic;
--    CLK_I7      : in  std_logic;
--    CLK_I8      : in  std_logic;

    PRE_SG_I    : in  std_logic;
    PRE_EN_I    : in  std_logic;

    PRE_IS_I1   : in  std_logic;
    PRE_IS_I2   : in  std_logic;
    PRE_IS_I3   : in  std_logic;
    PRE_IS_I4   : in  std_logic;

    MAIN_SG_I   : in  std_logic;

    MAIN_EN_I1  : in  std_logic;
    MAIN_EN_I2  : in  std_logic;
    MAIN_EN_I3  : in  std_logic;
    MAIN_EN_I4  : in  std_logic;
    MAIN_EN_I5  : in  std_logic;
    MAIN_EN_I6  : in  std_logic;

    MARG_S_I1   : in  std_logic;
    MARG_S_I2   : in  std_logic;
    MARG_S_I3   : in  std_logic;
    MARG_S_I4   : in  std_logic;

    MARG_IS_I1  : in  std_logic;
    MARG_IS_I2  : in  std_logic;
    MARG_IS_I3  : in  std_logic;
    MARG_IS_I4  : in  std_logic;

    MARG_SV_I1  : in  std_logic;
    MARG_SV_I2  : in  std_logic;
    MARG_SV_I3  : in  std_logic;
    MARG_SV_I4  : in  std_logic;
    MARG_SV_I5  : in  std_logic;

    MARG_ISV_I1 : in  std_logic;
    MARG_ISV_I2 : in  std_logic;
    MARG_ISV_I3 : in  std_logic;
    MARG_ISV_I4 : in  std_logic;
    MARG_ISV_I5 : in  std_logic;

    POST_EN_I1  : in  std_logic;
    POST_EN_I2  : in  std_logic;
    POST_EN_I3  : in  std_logic;
    POST_EN_I4  : in  std_logic;
    POST_EN_I5  : in  std_logic;

    POST_SG_I   : in  std_logic;

    POST_IS_I1  : in  std_logic;
    POST_IS_I2  : in  std_logic;
    POST_IS_I3  : in  std_logic;
    POST_IS_I4  : in  std_logic;

    POST_ISV_I1 : in  std_logic;
    POST_ISV_I2 : in  std_logic;
    POST_ISV_I3 : in  std_logic;
    POST_ISV_I4 : in  std_logic;

    TX_SEL_I1   : in  std_logic;
    TX_SEL_I2   : in  std_logic;
    TX_SEL_I3   : in  std_logic;
    TX_SEL_I4   : in  std_logic;
    TX_SEL_I5   : in  std_logic;
    TX_SEL_I6   : in  std_logic;

    CT_CAP_I1   : in  std_logic;
    CT_CAP_I2   : in  std_logic;
    CT_CAP_I3   : in  std_logic;
    CT_CAP_I4   : in  std_logic;

    CT_RESP_I1  : in  std_logic;
    CT_RESP_I2  : in  std_logic;
    CT_RESP_I3  : in  std_logic;
    CT_RESP_I4  : in  std_logic;

    CT_RESN_I1  : in  std_logic;
    CT_RESN_I2  : in  std_logic;
    CT_RESN_I3  : in  std_logic;
    CT_RESN_I4  : in  std_logic;

    M_EYE_I     : in  std_logic;

    RX_SEL_I1   : in  std_logic;
    RX_SEL_I2   : in  std_logic;
    RX_SEL_I3   : in  std_logic;
    RX_SEL_I4   : in  std_logic;
    RX_SEL_I5   : in  std_logic;
    RX_SEL_I6   : in  std_logic;

    PLL_RN_I    : in  std_logic;
    RST_N_I     : in  std_logic;

    CAL_1P_I1   : in  std_logic;
    CAL_1P_I2   : in  std_logic;
    CAL_1P_I3   : in  std_logic;
    CAL_1P_I4   : in  std_logic;
    CAL_1P_I5   : in  std_logic;
    CAL_1P_I6   : in  std_logic;
    CAL_1P_I7   : in  std_logic;
    CAL_1P_I8   : in  std_logic;

    CAL_2N_I1   : in  std_logic;
    CAL_2N_I2   : in  std_logic;
    CAL_2N_I3   : in  std_logic;
    CAL_2N_I4   : in  std_logic;
    CAL_2N_I5   : in  std_logic;
    CAL_2N_I6   : in  std_logic;
    CAL_2N_I7   : in  std_logic;
    CAL_2N_I8   : in  std_logic;

    CAL_3N_I1   : in  std_logic;
    CAL_3N_I2   : in  std_logic;
    CAL_3N_I3   : in  std_logic;
    CAL_3N_I4   : in  std_logic;
    CAL_3N_I5   : in  std_logic;
    CAL_3N_I6   : in  std_logic;
    CAL_3N_I7   : in  std_logic;
    CAL_3N_I8   : in  std_logic;

    CAL_4P_I1   : in  std_logic;
    CAL_4P_I2   : in  std_logic;
    CAL_4P_I3   : in  std_logic;
    CAL_4P_I4   : in  std_logic;
    CAL_4P_I5   : in  std_logic;
    CAL_4P_I6   : in  std_logic;
    CAL_4P_I7   : in  std_logic;
    CAL_4P_I8   : in  std_logic;

    CAL_SEL_I1  : in  std_logic;
    CAL_SEL_I2  : in  std_logic;
    CAL_SEL_I3  : in  std_logic;
    CAL_SEL_I4  : in  std_logic;

    CAL_E_I     : in  std_logic;
    LOCK_E_I    : in  std_logic;
    OVS_E_I     : in  std_logic;

    TST_I1      : in  std_logic;
    TST_I2      : in  std_logic;
    TST_I3      : in  std_logic;
    TST_I4      : in  std_logic;
    TST_I5      : in  std_logic;
    TST_I6      : in  std_logic;
    TST_I7      : in  std_logic;
    TST_I8      : in  std_logic;

    CLK_O       : out std_logic;
    LOCK_O      : out std_logic;
    CAL_O       : out std_logic;

    TST_O1      : out std_logic;
    TST_O2      : out std_logic;
    TST_O3      : out std_logic;
    TST_O4      : out std_logic;
    TST_O5      : out std_logic;
    TST_O6      : out std_logic;
    TST_O7      : out std_logic;
    TST_O8      : out std_logic;

    LINK_TX0    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX1    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX2    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX3    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX4    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX5    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_RX0    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX1    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX2    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX3    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX4    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX5    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);

    CLK_EXT_I   : in  std_logic
);
end component;
--#}}}#

begin

-- ctrl: NX_PMA_L#{{{#
ctrl: NX_PMA_L generic map (
    main_test                   => cfg_main_i(33 downto 26)
  , rx_pma_half_step            => cfg_main_i(25)
  , pll_pma_int_data_len        => cfg_main_i(24)
  , pll_pma_cpump_n             => cfg_main_i(23 downto 21)
  , pll_pma_divf                => cfg_main_i(20 downto 19)
  , pll_pma_divm                => cfg_main_i(18 downto 17)
  , pll_pma_divn                => cfg_main_i(16)
  , pll_pma_lvds_mux            => cfg_main_i(15)
  , pll_pma_mux_ckref           => cfg_main_i(14)
  , pll_pma_divf_en_n           => cfg_main_i(13)
  , pll_pma_divm_en_n           => cfg_main_i(12)
  , pll_pma_divn_en_n           => cfg_main_i(11)
  , main_clk_to_fabric_div_mode => cfg_main_i(10)
  , main_clk_to_fabric_div_en   => cfg_main_i(9)
  , main_clk_to_fabric_sel      => cfg_main_i(8)
  , main_use_only_usr_clock     => cfg_main_i(7)
  , main_use_pcs_clk_2          => cfg_main_i(6)
  , pcs_word_len                => cfg_main_i(5 downto 4)
  , pcs_ovs_mode                => cfg_main_i(3)
  , pcs_pll_lock_count          => cfg_main_i(2 downto 0)
  , location                    => location & ":COMMON1.PMA1"
 )
port map (
    CLK_USER_I  => hssl_clk_user_i
  , CLK_REF_I   => hssl_clk_ref_i
--    CLK_I1      => hssl_clock_i(0)
--  , CLK_I2      => hssl_clock_i(1)
--  , CLK_I3      => hssl_clock_i(2)
--  , CLK_I4      => hssl_clock_i(3)
--  , CLK_I5      => hssl_clock_i(4)
--  , CLK_I6      => hssl_clock_i(5)
--  , CLK_I7      => hssl_clock_i(6)
--  , CLK_I8      => hssl_clock_i(7)

  , PRE_SG_I    => usr_com_tx_pma_pre_sign_i
  , PRE_EN_I    => usr_com_tx_pma_pre_en_i

  , PRE_IS_I1   => usr_com_tx_pma_pre_input_sel_i(0)
  , PRE_IS_I2   => usr_com_tx_pma_pre_input_sel_i(1)
  , PRE_IS_I3   => usr_com_tx_pma_pre_input_sel_i(2)
  , PRE_IS_I4   => usr_com_tx_pma_pre_input_sel_i(3)

  , MAIN_SG_I   => usr_com_tx_pma_main_sign_i

  , MAIN_EN_I1  => usr_com_tx_pma_main_en_i(0)
  , MAIN_EN_I2  => usr_com_tx_pma_main_en_i(1)
  , MAIN_EN_I3  => usr_com_tx_pma_main_en_i(2)
  , MAIN_EN_I4  => usr_com_tx_pma_main_en_i(3)
  , MAIN_EN_I5  => usr_com_tx_pma_main_en_i(4)
  , MAIN_EN_I6  => usr_com_tx_pma_main_en_i(5)

  , MARG_S_I1   => usr_com_tx_pma_margin_sel_i(0)
  , MARG_S_I2   => usr_com_tx_pma_margin_sel_i(1)
  , MARG_S_I3   => usr_com_tx_pma_margin_sel_i(2)
  , MARG_S_I4   => usr_com_tx_pma_margin_sel_i(3)

  , MARG_IS_I1  => usr_com_tx_pma_margin_input_sel_i(0)
  , MARG_IS_I2  => usr_com_tx_pma_margin_input_sel_i(1)
  , MARG_IS_I3  => usr_com_tx_pma_margin_input_sel_i(2)
  , MARG_IS_I4  => usr_com_tx_pma_margin_input_sel_i(3)

  , MARG_SV_I1  => usr_com_tx_pma_margin_sel_var_i(0)
  , MARG_SV_I2  => usr_com_tx_pma_margin_sel_var_i(1)
  , MARG_SV_I3  => usr_com_tx_pma_margin_sel_var_i(2)
  , MARG_SV_I4  => usr_com_tx_pma_margin_sel_var_i(3)
  , MARG_SV_I5  => usr_com_tx_pma_margin_sel_var_i(4)

  , MARG_ISV_I1 => usr_com_tx_pma_margin_input_sel_var_i(0)
  , MARG_ISV_I2 => usr_com_tx_pma_margin_input_sel_var_i(1)
  , MARG_ISV_I3 => usr_com_tx_pma_margin_input_sel_var_i(2)
  , MARG_ISV_I4 => usr_com_tx_pma_margin_input_sel_var_i(3)
  , MARG_ISV_I5 => usr_com_tx_pma_margin_input_sel_var_i(4)

  , POST_EN_I1  => usr_com_tx_pma_post_en_i(0)
  , POST_EN_I2  => usr_com_tx_pma_post_en_i(1)
  , POST_EN_I3  => usr_com_tx_pma_post_en_i(2)
  , POST_EN_I4  => usr_com_tx_pma_post_en_i(3)
  , POST_EN_I5  => usr_com_tx_pma_post_en_i(4)

  , POST_SG_I   => usr_com_tx_pma_post_sign_i

  , POST_IS_I1  => usr_com_tx_pma_post_input_sel_i(0)
  , POST_IS_I2  => usr_com_tx_pma_post_input_sel_i(1)
  , POST_IS_I3  => usr_com_tx_pma_post_input_sel_i(2)
  , POST_IS_I4  => usr_com_tx_pma_post_input_sel_i(3)

  , POST_ISV_I1 => usr_com_tx_pma_post_input_sel_var_i(0)
  , POST_ISV_I2 => usr_com_tx_pma_post_input_sel_var_i(1)
  , POST_ISV_I3 => usr_com_tx_pma_post_input_sel_var_i(2)
  , POST_ISV_I4 => usr_com_tx_pma_post_input_sel_var_i(3)

  , TX_SEL_I1   => usr_com_ctrl_tx_sel_i(0)
  , TX_SEL_I2   => usr_com_ctrl_tx_sel_i(1)
  , TX_SEL_I3   => usr_com_ctrl_tx_sel_i(2)
  , TX_SEL_I4   => usr_com_ctrl_tx_sel_i(3)
  , TX_SEL_I5   => usr_com_ctrl_tx_sel_i(4)
  , TX_SEL_I6   => usr_com_ctrl_tx_sel_i(5)

  , CT_CAP_I1   => usr_com_rx_pma_ctle_cap_i(0)
  , CT_CAP_I2   => usr_com_rx_pma_ctle_cap_i(1)
  , CT_CAP_I3   => usr_com_rx_pma_ctle_cap_i(2)
  , CT_CAP_I4   => usr_com_rx_pma_ctle_cap_i(3)

  , CT_RESP_I1  => usr_com_rx_pma_ctle_resp_i(0)
  , CT_RESP_I2  => usr_com_rx_pma_ctle_resp_i(1)
  , CT_RESP_I3  => usr_com_rx_pma_ctle_resp_i(2)
  , CT_RESP_I4  => usr_com_rx_pma_ctle_resp_i(3)

  , CT_RESN_I1  => usr_com_rx_pma_ctle_resn_i(0)
  , CT_RESN_I2  => usr_com_rx_pma_ctle_resn_i(1)
  , CT_RESN_I3  => usr_com_rx_pma_ctle_resn_i(2)
  , CT_RESN_I4  => usr_com_rx_pma_ctle_resn_i(3)

  , M_EYE_I     => usr_com_rx_pma_m_eye_i

  , RX_SEL_I1   => usr_com_ctrl_rx_sel_i(0)
  , RX_SEL_I2   => usr_com_ctrl_rx_sel_i(1)
  , RX_SEL_I3   => usr_com_ctrl_rx_sel_i(2)
  , RX_SEL_I4   => usr_com_ctrl_rx_sel_i(3)
  , RX_SEL_I5   => usr_com_ctrl_rx_sel_i(4)
  , RX_SEL_I6   => usr_com_ctrl_rx_sel_i(5)

  , PLL_RN_I    => usr_pll_pma_rst_n_i
  , RST_N_I     => usr_main_rst_n_i

  , CAL_1P_I1   => usr_calibrate_pma_res_p1_i(0)
  , CAL_1P_I2   => usr_calibrate_pma_res_p1_i(1)
  , CAL_1P_I3   => usr_calibrate_pma_res_p1_i(2)
  , CAL_1P_I4   => usr_calibrate_pma_res_p1_i(3)
  , CAL_1P_I5   => usr_calibrate_pma_res_p1_i(4)
  , CAL_1P_I6   => usr_calibrate_pma_res_p1_i(5)
  , CAL_1P_I7   => usr_calibrate_pma_res_p1_i(6)
  , CAL_1P_I8   => usr_calibrate_pma_res_p1_i(7)

  , CAL_2N_I1   => usr_calibrate_pma_res_n2_i(0)
  , CAL_2N_I2   => usr_calibrate_pma_res_n2_i(1)
  , CAL_2N_I3   => usr_calibrate_pma_res_n2_i(2)
  , CAL_2N_I4   => usr_calibrate_pma_res_n2_i(3)
  , CAL_2N_I5   => usr_calibrate_pma_res_n2_i(4)
  , CAL_2N_I6   => usr_calibrate_pma_res_n2_i(5)
  , CAL_2N_I7   => usr_calibrate_pma_res_n2_i(6)
  , CAL_2N_I8   => usr_calibrate_pma_res_n2_i(7)

  , CAL_3N_I1   => usr_calibrate_pma_res_n3_i(0)
  , CAL_3N_I2   => usr_calibrate_pma_res_n3_i(1)
  , CAL_3N_I3   => usr_calibrate_pma_res_n3_i(2)
  , CAL_3N_I4   => usr_calibrate_pma_res_n3_i(3)
  , CAL_3N_I5   => usr_calibrate_pma_res_n3_i(4)
  , CAL_3N_I6   => usr_calibrate_pma_res_n3_i(5)
  , CAL_3N_I7   => usr_calibrate_pma_res_n3_i(6)
  , CAL_3N_I8   => usr_calibrate_pma_res_n3_i(7)

  , CAL_4P_I1   => usr_calibrate_pma_res_p4_i(0)
  , CAL_4P_I2   => usr_calibrate_pma_res_p4_i(1)
  , CAL_4P_I3   => usr_calibrate_pma_res_p4_i(2)
  , CAL_4P_I4   => usr_calibrate_pma_res_p4_i(3)
  , CAL_4P_I5   => usr_calibrate_pma_res_p4_i(4)
  , CAL_4P_I6   => usr_calibrate_pma_res_p4_i(5)
  , CAL_4P_I7   => usr_calibrate_pma_res_p4_i(6)
  , CAL_4P_I8   => usr_calibrate_pma_res_p4_i(7)

  , CAL_SEL_I1  => usr_calibrate_pma_sel_i(0)
  , CAL_SEL_I2  => usr_calibrate_pma_sel_i(1)
  , CAL_SEL_I3  => usr_calibrate_pma_sel_i(2)
  , CAL_SEL_I4  => usr_calibrate_pma_sel_i(3)

  , CAL_E_I     => usr_calibrate_pma_en_i
  , LOCK_E_I    => usr_pcs_ctrl_pll_lock_en_i
  , OVS_E_I     => usr_pcs_ctrl_ovs_en_i

  , TST_I1      => usr_main_test_i(0)
  , TST_I2      => usr_main_test_i(1)
  , TST_I3      => usr_main_test_i(2)
  , TST_I4      => usr_main_test_i(3)
  , TST_I5      => usr_main_test_i(4)
  , TST_I6      => usr_main_test_i(5)
  , TST_I7      => usr_main_test_i(6)
  , TST_I8      => usr_main_test_i(7)

  , CLK_O       => hssl_clock_o
  , LOCK_O      => usr_pll_lock_o
  , CAL_O       => usr_calibrate_pma_out_o

  , TST_O1      => usr_main_test_o(0)
  , TST_O2      => usr_main_test_o(1)
  , TST_O3      => usr_main_test_o(2)
  , TST_O4      => usr_main_test_o(3)
  , TST_O5      => usr_main_test_o(4)
  , TST_O6      => usr_main_test_o(5)
  , TST_O7      => usr_main_test_o(6)
  , TST_O8      => usr_main_test_o(7)

  , LINK_TX0    => LINK_TX0
  , LINK_TX1    => LINK_TX1
  , LINK_TX2    => LINK_TX2
  , LINK_TX3    => LINK_TX3
  , LINK_TX4    => LINK_TX4
  , LINK_TX5    => LINK_TX5
  , LINK_RX0    => LINK_RX0
  , LINK_RX1    => LINK_RX1
  , LINK_RX2    => LINK_RX2
  , LINK_RX3    => LINK_RX3
  , LINK_RX4    => LINK_RX4
  , LINK_RX5    => LINK_RX5

  , CLK_EXT_I   => pma_clk_ext_i
);
--#}}}#

-- txlane0: NX_CTX_L#{{{#
txlane0: NX_CTX_L generic map (
   pma_clk_pos          => cfg_tx0_i(31)
 , pcs_protocol_size    => cfg_tx0_i(30)
 , pcs_8b_scr_sel       => cfg_tx0_i(29)
 , pcs_scr_init         => cfg_tx0_i(28 downto 12)
 , pcs_scr_bypass       => cfg_tx0_i(11)
 , pcs_sync_supported   => cfg_tx0_i(10)
 , pcs_replace_bypass   => cfg_tx0_i(9)
 , pcs_enc_bypass       => cfg_tx0_i(8)
 , pcs_loopback         => cfg_tx0_i(7)
 , pcs_polarity         => cfg_tx0_i(6)
 , pcs_esistream_fsm_en => cfg_tx0_i(5)
 , test                 => cfg_tx0_i(4 downto 3)
 , pcs_bypass_pma_cdc   => cfg_tx0_i(2)
 , pcs_bypass_usr_cdc   => cfg_tx0_i(1)
 , pma_loopback         => cfg_tx0_i(0)
 , location             => location & ":CHANNEL1.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx0_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx0_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx0_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx0_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx0_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx0_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx0_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx0_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx0_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx0_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx0_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx0_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx0_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx0_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx0_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx0_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx0_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx0_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx0_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx0_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx0_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx0_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx0_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx0_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx0_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx0_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx0_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx0_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx0_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx0_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx0_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx0_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx0_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx0_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx0_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx0_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx0_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx0_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx0_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx0_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx0_ctrl_replace_en_i
  , RST_N_I  => usr_tx0_rst_n_i

  , TST_I1   => usr_tx0_test_i(0)
  , TST_I2   => usr_tx0_test_i(1)
  , TST_I3   => usr_tx0_test_i(2)
  , TST_I4   => usr_tx0_test_i(3)

  , DATA_I1  => usr_tx0_data_i(0)
  , DATA_I2  => usr_tx0_data_i(1)
  , DATA_I3  => usr_tx0_data_i(2)
  , DATA_I4  => usr_tx0_data_i(3)
  , DATA_I5  => usr_tx0_data_i(4)
  , DATA_I6  => usr_tx0_data_i(5)
  , DATA_I7  => usr_tx0_data_i(6)
  , DATA_I8  => usr_tx0_data_i(7)
  , DATA_I9  => usr_tx0_data_i(8)
  , DATA_I10 => usr_tx0_data_i(9)
  , DATA_I11 => usr_tx0_data_i(10)
  , DATA_I12 => usr_tx0_data_i(11)
  , DATA_I13 => usr_tx0_data_i(12)
  , DATA_I14 => usr_tx0_data_i(13)
  , DATA_I15 => usr_tx0_data_i(14)
  , DATA_I16 => usr_tx0_data_i(15)
  , DATA_I17 => usr_tx0_data_i(16)
  , DATA_I18 => usr_tx0_data_i(17)
  , DATA_I19 => usr_tx0_data_i(18)
  , DATA_I20 => usr_tx0_data_i(19)
  , DATA_I21 => usr_tx0_data_i(20)
  , DATA_I22 => usr_tx0_data_i(21)
  , DATA_I23 => usr_tx0_data_i(22)
  , DATA_I24 => usr_tx0_data_i(23)
  , DATA_I25 => usr_tx0_data_i(24)
  , DATA_I26 => usr_tx0_data_i(25)
  , DATA_I27 => usr_tx0_data_i(26)
  , DATA_I28 => usr_tx0_data_i(27)
  , DATA_I29 => usr_tx0_data_i(28)
  , DATA_I30 => usr_tx0_data_i(29)
  , DATA_I31 => usr_tx0_data_i(30)
  , DATA_I32 => usr_tx0_data_i(31)
  , DATA_I33 => usr_tx0_data_i(32)
  , DATA_I34 => usr_tx0_data_i(33)
  , DATA_I35 => usr_tx0_data_i(34)
  , DATA_I36 => usr_tx0_data_i(35)
  , DATA_I37 => usr_tx0_data_i(36)
  , DATA_I38 => usr_tx0_data_i(37)
  , DATA_I39 => usr_tx0_data_i(38)
  , DATA_I40 => usr_tx0_data_i(39)
  , DATA_I41 => usr_tx0_data_i(40)
  , DATA_I42 => usr_tx0_data_i(41)
  , DATA_I43 => usr_tx0_data_i(42)
  , DATA_I44 => usr_tx0_data_i(43)
  , DATA_I45 => usr_tx0_data_i(44)
  , DATA_I46 => usr_tx0_data_i(45)
  , DATA_I47 => usr_tx0_data_i(46)
  , DATA_I48 => usr_tx0_data_i(47)
  , DATA_I49 => usr_tx0_data_i(48)
  , DATA_I50 => usr_tx0_data_i(49)
  , DATA_I51 => usr_tx0_data_i(50)
  , DATA_I52 => usr_tx0_data_i(51)
  , DATA_I53 => usr_tx0_data_i(52)
  , DATA_I54 => usr_tx0_data_i(53)
  , DATA_I55 => usr_tx0_data_i(54)
  , DATA_I56 => usr_tx0_data_i(55)
  , DATA_I57 => usr_tx0_data_i(56)
  , DATA_I58 => usr_tx0_data_i(57)
  , DATA_I59 => usr_tx0_data_i(58)
  , DATA_I60 => usr_tx0_data_i(59)
  , DATA_I61 => usr_tx0_data_i(60)
  , DATA_I62 => usr_tx0_data_i(61)
  , DATA_I63 => usr_tx0_data_i(62)
  , DATA_I64 => usr_tx0_data_i(63)

  , TST_O1   => usr_tx0_test_o(0)
  , TST_O2   => usr_tx0_test_o(1)
  , TST_O3   => usr_tx0_test_o(2)
  , TST_O4   => usr_tx0_test_o(3)

  , BUSY_O   => usr_tx0_busy_o
  , CLK_E_I  => usr_tx0_pma_clk_en_i

  , LINK     => LINK_TX0

  , TX_O     => pma_tx0_o
);
--#}}}#

-- rxlane0: NX_CRX_L#{{{#
rxlane0: NX_CRX_L generic map (
    test                         => cfg_rx0_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx0_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx0_i(156)
  , pcs_debug_en                 => cfg_rx0_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx0_i(154)
  , pma_clk_pos                  => cfg_rx0_i(153)
  , pcs_protocol_size            => cfg_rx0_i(152)
  , pcs_loopback                 => cfg_rx0_i(151)
  , pcs_polarity                 => cfg_rx0_i(150)
  , pcs_p_comma_en               => cfg_rx0_i(149)
  , pcs_p_comma_val              => cfg_rx0_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx0_i(138)
  , pcs_m_comma_val              => cfg_rx0_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx0_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx0_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx0_i(115)
  , pcs_dec_bypass               => cfg_rx0_i(114)
  , pcs_el_buff_max_comp         => cfg_rx0_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx0_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx0_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx0_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx0_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx0_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx0_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx0_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx0_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx0_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx0_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx0_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx0_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx0_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx0_i(29)
  , pcs_buffers_bypass           => cfg_rx0_i(28)
  , pcs_sync_supported           => cfg_rx0_i(27)
  , pcs_replace_bypass           => cfg_rx0_i(26)
  , pcs_dscr_bypass              => cfg_rx0_i(25)
  , pcs_8b_dscr_sel              => cfg_rx0_i(24)
  , pcs_fsm_sel                  => cfg_rx0_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx0_i(21)
  , pma_pll_divm_en_n            => cfg_rx0_i(20)
  , pma_pll_divn_en_n            => cfg_rx0_i(19)
  , pma_cdr_cp                   => cfg_rx0_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx0_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx0_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx0_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx0_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx0_i(1)
  , pma_loopback                 => cfg_rx0_i(0)
  , location                     => location & ":CHANNEL1.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx0_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx0_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx0_ctrl_align_en_i
  , ALIGN_S_I => usr_rx0_ctrl_align_sync_i
  , REP_E_I   => usr_rx0_ctrl_replace_en_i
  , BUF_R_I   => usr_rx0_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx0_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx0_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx0_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx0_rst_n_i
  , CDR_R_I   => usr_rx0_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx0_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx0_pma_pll_rst_n_i

  , TST_I1    => usr_rx0_test_i(0)
  , TST_I2    => usr_rx0_test_i(1)
  , TST_I3    => usr_rx0_test_i(2)
  , TST_I4    => usr_rx0_test_i(3)

  , LOS_O     => usr_rx0_pma_loss_of_signal_o

  , DATA_O1   => usr_rx0_data_o(0)
  , DATA_O2   => usr_rx0_data_o(1)
  , DATA_O3   => usr_rx0_data_o(2)
  , DATA_O4   => usr_rx0_data_o(3)
  , DATA_O5   => usr_rx0_data_o(4)
  , DATA_O6   => usr_rx0_data_o(5)
  , DATA_O7   => usr_rx0_data_o(6)
  , DATA_O8   => usr_rx0_data_o(7)
  , DATA_O9   => usr_rx0_data_o(8)
  , DATA_O10  => usr_rx0_data_o(9)
  , DATA_O11  => usr_rx0_data_o(10)
  , DATA_O12  => usr_rx0_data_o(11)
  , DATA_O13  => usr_rx0_data_o(12)
  , DATA_O14  => usr_rx0_data_o(13)
  , DATA_O15  => usr_rx0_data_o(14)
  , DATA_O16  => usr_rx0_data_o(15)
  , DATA_O17  => usr_rx0_data_o(16)
  , DATA_O18  => usr_rx0_data_o(17)
  , DATA_O19  => usr_rx0_data_o(18)
  , DATA_O20  => usr_rx0_data_o(19)
  , DATA_O21  => usr_rx0_data_o(20)
  , DATA_O22  => usr_rx0_data_o(21)
  , DATA_O23  => usr_rx0_data_o(22)
  , DATA_O24  => usr_rx0_data_o(23)
  , DATA_O25  => usr_rx0_data_o(24)
  , DATA_O26  => usr_rx0_data_o(25)
  , DATA_O27  => usr_rx0_data_o(26)
  , DATA_O28  => usr_rx0_data_o(27)
  , DATA_O29  => usr_rx0_data_o(28)
  , DATA_O30  => usr_rx0_data_o(29)
  , DATA_O31  => usr_rx0_data_o(30)
  , DATA_O32  => usr_rx0_data_o(31)
  , DATA_O33  => usr_rx0_data_o(32)
  , DATA_O34  => usr_rx0_data_o(33)
  , DATA_O35  => usr_rx0_data_o(34)
  , DATA_O36  => usr_rx0_data_o(35)
  , DATA_O37  => usr_rx0_data_o(36)
  , DATA_O38  => usr_rx0_data_o(37)
  , DATA_O39  => usr_rx0_data_o(38)
  , DATA_O40  => usr_rx0_data_o(39)
  , DATA_O41  => usr_rx0_data_o(40)
  , DATA_O42  => usr_rx0_data_o(41)
  , DATA_O43  => usr_rx0_data_o(42)
  , DATA_O44  => usr_rx0_data_o(43)
  , DATA_O45  => usr_rx0_data_o(44)
  , DATA_O46  => usr_rx0_data_o(45)
  , DATA_O47  => usr_rx0_data_o(46)
  , DATA_O48  => usr_rx0_data_o(47)
  , DATA_O49  => usr_rx0_data_o(48)
  , DATA_O50  => usr_rx0_data_o(49)
  , DATA_O51  => usr_rx0_data_o(50)
  , DATA_O52  => usr_rx0_data_o(51)
  , DATA_O53  => usr_rx0_data_o(52)
  , DATA_O54  => usr_rx0_data_o(53)
  , DATA_O55  => usr_rx0_data_o(54)
  , DATA_O56  => usr_rx0_data_o(55)
  , DATA_O57  => usr_rx0_data_o(56)
  , DATA_O58  => usr_rx0_data_o(57)
  , DATA_O59  => usr_rx0_data_o(58)
  , DATA_O60  => usr_rx0_data_o(59)
  , DATA_O61  => usr_rx0_data_o(60)
  , DATA_O62  => usr_rx0_data_o(61)
  , DATA_O63  => usr_rx0_data_o(62)
  , DATA_O64  => usr_rx0_data_o(63)

  , CH_COM_O1 => usr_rx0_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx0_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx0_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx0_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx0_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx0_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx0_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx0_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx0_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx0_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx0_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx0_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx0_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx0_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx0_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx0_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx0_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx0_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx0_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx0_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx0_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx0_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx0_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx0_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx0_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx0_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx0_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx0_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx0_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx0_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx0_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx0_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx0_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx0_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx0_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx0_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx0_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx0_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx0_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx0_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx0_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx0_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx0_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx0_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx0_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx0_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx0_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx0_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx0_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx0_busy_o

  , TST_O1    => usr_rx0_test_o(0)
  , TST_O2    => usr_rx0_test_o(1)
  , TST_O3    => usr_rx0_test_o(2)
  , TST_O4    => usr_rx0_test_o(3)
  , TST_O5    => usr_rx0_test_o(4)
  , TST_O6    => usr_rx0_test_o(5)
  , TST_O7    => usr_rx0_test_o(6)
  , TST_O8    => usr_rx0_test_o(7)

  , LOCK_O    => usr_rx0_pll_lock_o

  , LINK      => LINK_RX0

  , RX_I      => pma_rx0_i
);
--#}}}#

-- txlane1: NX_CTX_L#{{{#
txlane1: NX_CTX_L generic map (
   pma_clk_pos          => cfg_tx1_i(31)
 , pcs_protocol_size    => cfg_tx1_i(30)
 , pcs_8b_scr_sel       => cfg_tx1_i(29)
 , pcs_scr_init         => cfg_tx1_i(28 downto 12)
 , pcs_scr_bypass       => cfg_tx1_i(11)
 , pcs_sync_supported   => cfg_tx1_i(10)
 , pcs_replace_bypass   => cfg_tx1_i(9)
 , pcs_enc_bypass       => cfg_tx1_i(8)
 , pcs_loopback         => cfg_tx1_i(7)
 , pcs_polarity         => cfg_tx1_i(6)
 , pcs_esistream_fsm_en => cfg_tx1_i(5)
 , test                 => cfg_tx1_i(4 downto 3)
 , pcs_bypass_pma_cdc   => cfg_tx1_i(2)
 , pcs_bypass_usr_cdc   => cfg_tx1_i(1)
 , pma_loopback         => cfg_tx1_i(0)
 , location             => location & ":CHANNEL2.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx1_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx1_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx1_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx1_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx1_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx1_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx1_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx1_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx1_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx1_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx1_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx1_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx1_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx1_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx1_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx1_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx1_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx1_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx1_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx1_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx1_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx1_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx1_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx1_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx1_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx1_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx1_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx1_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx1_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx1_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx1_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx1_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx1_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx1_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx1_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx1_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx1_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx1_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx1_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx1_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx1_ctrl_replace_en_i
  , RST_N_I  => usr_tx1_rst_n_i

  , TST_I1   => usr_tx1_test_i(0)
  , TST_I2   => usr_tx1_test_i(1)
  , TST_I3   => usr_tx1_test_i(2)
  , TST_I4   => usr_tx1_test_i(3)

  , DATA_I1  => usr_tx1_data_i(0)
  , DATA_I2  => usr_tx1_data_i(1)
  , DATA_I3  => usr_tx1_data_i(2)
  , DATA_I4  => usr_tx1_data_i(3)
  , DATA_I5  => usr_tx1_data_i(4)
  , DATA_I6  => usr_tx1_data_i(5)
  , DATA_I7  => usr_tx1_data_i(6)
  , DATA_I8  => usr_tx1_data_i(7)
  , DATA_I9  => usr_tx1_data_i(8)
  , DATA_I10 => usr_tx1_data_i(9)
  , DATA_I11 => usr_tx1_data_i(10)
  , DATA_I12 => usr_tx1_data_i(11)
  , DATA_I13 => usr_tx1_data_i(12)
  , DATA_I14 => usr_tx1_data_i(13)
  , DATA_I15 => usr_tx1_data_i(14)
  , DATA_I16 => usr_tx1_data_i(15)
  , DATA_I17 => usr_tx1_data_i(16)
  , DATA_I18 => usr_tx1_data_i(17)
  , DATA_I19 => usr_tx1_data_i(18)
  , DATA_I20 => usr_tx1_data_i(19)
  , DATA_I21 => usr_tx1_data_i(20)
  , DATA_I22 => usr_tx1_data_i(21)
  , DATA_I23 => usr_tx1_data_i(22)
  , DATA_I24 => usr_tx1_data_i(23)
  , DATA_I25 => usr_tx1_data_i(24)
  , DATA_I26 => usr_tx1_data_i(25)
  , DATA_I27 => usr_tx1_data_i(26)
  , DATA_I28 => usr_tx1_data_i(27)
  , DATA_I29 => usr_tx1_data_i(28)
  , DATA_I30 => usr_tx1_data_i(29)
  , DATA_I31 => usr_tx1_data_i(30)
  , DATA_I32 => usr_tx1_data_i(31)
  , DATA_I33 => usr_tx1_data_i(32)
  , DATA_I34 => usr_tx1_data_i(33)
  , DATA_I35 => usr_tx1_data_i(34)
  , DATA_I36 => usr_tx1_data_i(35)
  , DATA_I37 => usr_tx1_data_i(36)
  , DATA_I38 => usr_tx1_data_i(37)
  , DATA_I39 => usr_tx1_data_i(38)
  , DATA_I40 => usr_tx1_data_i(39)
  , DATA_I41 => usr_tx1_data_i(40)
  , DATA_I42 => usr_tx1_data_i(41)
  , DATA_I43 => usr_tx1_data_i(42)
  , DATA_I44 => usr_tx1_data_i(43)
  , DATA_I45 => usr_tx1_data_i(44)
  , DATA_I46 => usr_tx1_data_i(45)
  , DATA_I47 => usr_tx1_data_i(46)
  , DATA_I48 => usr_tx1_data_i(47)
  , DATA_I49 => usr_tx1_data_i(48)
  , DATA_I50 => usr_tx1_data_i(49)
  , DATA_I51 => usr_tx1_data_i(50)
  , DATA_I52 => usr_tx1_data_i(51)
  , DATA_I53 => usr_tx1_data_i(52)
  , DATA_I54 => usr_tx1_data_i(53)
  , DATA_I55 => usr_tx1_data_i(54)
  , DATA_I56 => usr_tx1_data_i(55)
  , DATA_I57 => usr_tx1_data_i(56)
  , DATA_I58 => usr_tx1_data_i(57)
  , DATA_I59 => usr_tx1_data_i(58)
  , DATA_I60 => usr_tx1_data_i(59)
  , DATA_I61 => usr_tx1_data_i(60)
  , DATA_I62 => usr_tx1_data_i(61)
  , DATA_I63 => usr_tx1_data_i(62)
  , DATA_I64 => usr_tx1_data_i(63)

  , TST_O1   => usr_tx1_test_o(0)
  , TST_O2   => usr_tx1_test_o(1)
  , TST_O3   => usr_tx1_test_o(2)
  , TST_O4   => usr_tx1_test_o(3)

  , BUSY_O   => usr_tx1_busy_o
  , CLK_E_I  => usr_tx1_pma_clk_en_i

  , LINK     => LINK_TX1

  , TX_O     => pma_tx1_o
);
--#}}}#

-- rxlane1: NX_CRX_L#{{{#
rxlane1: NX_CRX_L generic map (
    test                         => cfg_rx1_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx1_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx1_i(156)
  , pcs_debug_en                 => cfg_rx1_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx1_i(154)
  , pma_clk_pos                  => cfg_rx1_i(153)
  , pcs_protocol_size            => cfg_rx1_i(152)
  , pcs_loopback                 => cfg_rx1_i(151)
  , pcs_polarity                 => cfg_rx1_i(150)
  , pcs_p_comma_en               => cfg_rx1_i(149)
  , pcs_p_comma_val              => cfg_rx1_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx1_i(138)
  , pcs_m_comma_val              => cfg_rx1_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx1_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx1_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx1_i(115)
  , pcs_dec_bypass               => cfg_rx1_i(114)
  , pcs_el_buff_max_comp         => cfg_rx1_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx1_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx1_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx1_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx1_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx1_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx1_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx1_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx1_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx1_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx1_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx1_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx1_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx1_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx1_i(29)
  , pcs_buffers_bypass           => cfg_rx1_i(28)
  , pcs_sync_supported           => cfg_rx1_i(27)
  , pcs_replace_bypass           => cfg_rx1_i(26)
  , pcs_dscr_bypass              => cfg_rx1_i(25)
  , pcs_8b_dscr_sel              => cfg_rx1_i(24)
  , pcs_fsm_sel                  => cfg_rx1_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx1_i(21)
  , pma_pll_divm_en_n            => cfg_rx1_i(20)
  , pma_pll_divn_en_n            => cfg_rx1_i(19)
  , pma_cdr_cp                   => cfg_rx1_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx1_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx1_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx1_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx1_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx1_i(1)
  , pma_loopback                 => cfg_rx1_i(0)
  , location                     => location & ":CHANNEL2.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx1_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx1_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx1_ctrl_align_en_i
  , ALIGN_S_I => usr_rx1_ctrl_align_sync_i
  , REP_E_I   => usr_rx1_ctrl_replace_en_i
  , BUF_R_I   => usr_rx1_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx1_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx1_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx1_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx1_rst_n_i
  , CDR_R_I   => usr_rx1_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx1_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx1_pma_pll_rst_n_i

  , TST_I1    => usr_rx1_test_i(0)
  , TST_I2    => usr_rx1_test_i(1)
  , TST_I3    => usr_rx1_test_i(2)
  , TST_I4    => usr_rx1_test_i(3)

  , LOS_O     => usr_rx1_pma_loss_of_signal_o

  , DATA_O1   => usr_rx1_data_o(0)
  , DATA_O2   => usr_rx1_data_o(1)
  , DATA_O3   => usr_rx1_data_o(2)
  , DATA_O4   => usr_rx1_data_o(3)
  , DATA_O5   => usr_rx1_data_o(4)
  , DATA_O6   => usr_rx1_data_o(5)
  , DATA_O7   => usr_rx1_data_o(6)
  , DATA_O8   => usr_rx1_data_o(7)
  , DATA_O9   => usr_rx1_data_o(8)
  , DATA_O10  => usr_rx1_data_o(9)
  , DATA_O11  => usr_rx1_data_o(10)
  , DATA_O12  => usr_rx1_data_o(11)
  , DATA_O13  => usr_rx1_data_o(12)
  , DATA_O14  => usr_rx1_data_o(13)
  , DATA_O15  => usr_rx1_data_o(14)
  , DATA_O16  => usr_rx1_data_o(15)
  , DATA_O17  => usr_rx1_data_o(16)
  , DATA_O18  => usr_rx1_data_o(17)
  , DATA_O19  => usr_rx1_data_o(18)
  , DATA_O20  => usr_rx1_data_o(19)
  , DATA_O21  => usr_rx1_data_o(20)
  , DATA_O22  => usr_rx1_data_o(21)
  , DATA_O23  => usr_rx1_data_o(22)
  , DATA_O24  => usr_rx1_data_o(23)
  , DATA_O25  => usr_rx1_data_o(24)
  , DATA_O26  => usr_rx1_data_o(25)
  , DATA_O27  => usr_rx1_data_o(26)
  , DATA_O28  => usr_rx1_data_o(27)
  , DATA_O29  => usr_rx1_data_o(28)
  , DATA_O30  => usr_rx1_data_o(29)
  , DATA_O31  => usr_rx1_data_o(30)
  , DATA_O32  => usr_rx1_data_o(31)
  , DATA_O33  => usr_rx1_data_o(32)
  , DATA_O34  => usr_rx1_data_o(33)
  , DATA_O35  => usr_rx1_data_o(34)
  , DATA_O36  => usr_rx1_data_o(35)
  , DATA_O37  => usr_rx1_data_o(36)
  , DATA_O38  => usr_rx1_data_o(37)
  , DATA_O39  => usr_rx1_data_o(38)
  , DATA_O40  => usr_rx1_data_o(39)
  , DATA_O41  => usr_rx1_data_o(40)
  , DATA_O42  => usr_rx1_data_o(41)
  , DATA_O43  => usr_rx1_data_o(42)
  , DATA_O44  => usr_rx1_data_o(43)
  , DATA_O45  => usr_rx1_data_o(44)
  , DATA_O46  => usr_rx1_data_o(45)
  , DATA_O47  => usr_rx1_data_o(46)
  , DATA_O48  => usr_rx1_data_o(47)
  , DATA_O49  => usr_rx1_data_o(48)
  , DATA_O50  => usr_rx1_data_o(49)
  , DATA_O51  => usr_rx1_data_o(50)
  , DATA_O52  => usr_rx1_data_o(51)
  , DATA_O53  => usr_rx1_data_o(52)
  , DATA_O54  => usr_rx1_data_o(53)
  , DATA_O55  => usr_rx1_data_o(54)
  , DATA_O56  => usr_rx1_data_o(55)
  , DATA_O57  => usr_rx1_data_o(56)
  , DATA_O58  => usr_rx1_data_o(57)
  , DATA_O59  => usr_rx1_data_o(58)
  , DATA_O60  => usr_rx1_data_o(59)
  , DATA_O61  => usr_rx1_data_o(60)
  , DATA_O62  => usr_rx1_data_o(61)
  , DATA_O63  => usr_rx1_data_o(62)
  , DATA_O64  => usr_rx1_data_o(63)

  , CH_COM_O1 => usr_rx1_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx1_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx1_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx1_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx1_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx1_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx1_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx1_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx1_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx1_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx1_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx1_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx1_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx1_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx1_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx1_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx1_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx1_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx1_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx1_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx1_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx1_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx1_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx1_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx1_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx1_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx1_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx1_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx1_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx1_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx1_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx1_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx1_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx1_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx1_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx1_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx1_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx1_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx1_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx1_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx1_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx1_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx1_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx1_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx1_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx1_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx1_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx1_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx1_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx1_busy_o

  , TST_O1    => usr_rx1_test_o(0)
  , TST_O2    => usr_rx1_test_o(1)
  , TST_O3    => usr_rx1_test_o(2)
  , TST_O4    => usr_rx1_test_o(3)
  , TST_O5    => usr_rx1_test_o(4)
  , TST_O6    => usr_rx1_test_o(5)
  , TST_O7    => usr_rx1_test_o(6)
  , TST_O8    => usr_rx1_test_o(7)

  , LOCK_O    => usr_rx1_pll_lock_o

  , LINK      => LINK_RX1

  , RX_I      => pma_rx1_i
);
--#}}}#

-- txlane2: NX_CTX_L#{{{#
txlane2: NX_CTX_L generic map (
   pma_clk_pos          => cfg_tx2_i(31)
 , pcs_protocol_size    => cfg_tx2_i(30)
 , pcs_8b_scr_sel       => cfg_tx2_i(29)
 , pcs_scr_init         => cfg_tx2_i(28 downto 12)
 , pcs_scr_bypass       => cfg_tx2_i(11)
 , pcs_sync_supported   => cfg_tx2_i(10)
 , pcs_replace_bypass   => cfg_tx2_i(9)
 , pcs_enc_bypass       => cfg_tx2_i(8)
 , pcs_loopback         => cfg_tx2_i(7)
 , pcs_polarity         => cfg_tx2_i(6)
 , pcs_esistream_fsm_en => cfg_tx2_i(5)
 , test                 => cfg_tx2_i(4 downto 3)
 , pcs_bypass_pma_cdc   => cfg_tx2_i(2)
 , pcs_bypass_usr_cdc   => cfg_tx2_i(1)
 , pma_loopback         => cfg_tx2_i(0)
 , location             => location & ":CHANNEL3.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx2_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx2_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx2_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx2_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx2_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx2_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx2_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx2_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx2_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx2_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx2_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx2_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx2_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx2_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx2_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx2_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx2_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx2_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx2_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx2_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx2_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx2_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx2_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx2_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx2_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx2_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx2_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx2_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx2_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx2_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx2_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx2_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx2_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx2_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx2_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx2_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx2_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx2_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx2_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx2_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx2_ctrl_replace_en_i
  , RST_N_I  => usr_tx2_rst_n_i

  , TST_I1   => usr_tx2_test_i(0)
  , TST_I2   => usr_tx2_test_i(1)
  , TST_I3   => usr_tx2_test_i(2)
  , TST_I4   => usr_tx2_test_i(3)

  , DATA_I1  => usr_tx2_data_i(0)
  , DATA_I2  => usr_tx2_data_i(1)
  , DATA_I3  => usr_tx2_data_i(2)
  , DATA_I4  => usr_tx2_data_i(3)
  , DATA_I5  => usr_tx2_data_i(4)
  , DATA_I6  => usr_tx2_data_i(5)
  , DATA_I7  => usr_tx2_data_i(6)
  , DATA_I8  => usr_tx2_data_i(7)
  , DATA_I9  => usr_tx2_data_i(8)
  , DATA_I10 => usr_tx2_data_i(9)
  , DATA_I11 => usr_tx2_data_i(10)
  , DATA_I12 => usr_tx2_data_i(11)
  , DATA_I13 => usr_tx2_data_i(12)
  , DATA_I14 => usr_tx2_data_i(13)
  , DATA_I15 => usr_tx2_data_i(14)
  , DATA_I16 => usr_tx2_data_i(15)
  , DATA_I17 => usr_tx2_data_i(16)
  , DATA_I18 => usr_tx2_data_i(17)
  , DATA_I19 => usr_tx2_data_i(18)
  , DATA_I20 => usr_tx2_data_i(19)
  , DATA_I21 => usr_tx2_data_i(20)
  , DATA_I22 => usr_tx2_data_i(21)
  , DATA_I23 => usr_tx2_data_i(22)
  , DATA_I24 => usr_tx2_data_i(23)
  , DATA_I25 => usr_tx2_data_i(24)
  , DATA_I26 => usr_tx2_data_i(25)
  , DATA_I27 => usr_tx2_data_i(26)
  , DATA_I28 => usr_tx2_data_i(27)
  , DATA_I29 => usr_tx2_data_i(28)
  , DATA_I30 => usr_tx2_data_i(29)
  , DATA_I31 => usr_tx2_data_i(30)
  , DATA_I32 => usr_tx2_data_i(31)
  , DATA_I33 => usr_tx2_data_i(32)
  , DATA_I34 => usr_tx2_data_i(33)
  , DATA_I35 => usr_tx2_data_i(34)
  , DATA_I36 => usr_tx2_data_i(35)
  , DATA_I37 => usr_tx2_data_i(36)
  , DATA_I38 => usr_tx2_data_i(37)
  , DATA_I39 => usr_tx2_data_i(38)
  , DATA_I40 => usr_tx2_data_i(39)
  , DATA_I41 => usr_tx2_data_i(40)
  , DATA_I42 => usr_tx2_data_i(41)
  , DATA_I43 => usr_tx2_data_i(42)
  , DATA_I44 => usr_tx2_data_i(43)
  , DATA_I45 => usr_tx2_data_i(44)
  , DATA_I46 => usr_tx2_data_i(45)
  , DATA_I47 => usr_tx2_data_i(46)
  , DATA_I48 => usr_tx2_data_i(47)
  , DATA_I49 => usr_tx2_data_i(48)
  , DATA_I50 => usr_tx2_data_i(49)
  , DATA_I51 => usr_tx2_data_i(50)
  , DATA_I52 => usr_tx2_data_i(51)
  , DATA_I53 => usr_tx2_data_i(52)
  , DATA_I54 => usr_tx2_data_i(53)
  , DATA_I55 => usr_tx2_data_i(54)
  , DATA_I56 => usr_tx2_data_i(55)
  , DATA_I57 => usr_tx2_data_i(56)
  , DATA_I58 => usr_tx2_data_i(57)
  , DATA_I59 => usr_tx2_data_i(58)
  , DATA_I60 => usr_tx2_data_i(59)
  , DATA_I61 => usr_tx2_data_i(60)
  , DATA_I62 => usr_tx2_data_i(61)
  , DATA_I63 => usr_tx2_data_i(62)
  , DATA_I64 => usr_tx2_data_i(63)

  , TST_O1   => usr_tx2_test_o(0)
  , TST_O2   => usr_tx2_test_o(1)
  , TST_O3   => usr_tx2_test_o(2)
  , TST_O4   => usr_tx2_test_o(3)

  , BUSY_O   => usr_tx2_busy_o
  , CLK_E_I  => usr_tx2_pma_clk_en_i

  , LINK     => LINK_TX2

  , TX_O     => pma_tx2_o
);
--#}}}#

-- rxlane2: NX_CRX_L#{{{#
rxlane2: NX_CRX_L generic map (
    test                         => cfg_rx2_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx2_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx2_i(156)
  , pcs_debug_en                 => cfg_rx2_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx2_i(154)
  , pma_clk_pos                  => cfg_rx2_i(153)
  , pcs_protocol_size            => cfg_rx2_i(152)
  , pcs_loopback                 => cfg_rx2_i(151)
  , pcs_polarity                 => cfg_rx2_i(150)
  , pcs_p_comma_en               => cfg_rx2_i(149)
  , pcs_p_comma_val              => cfg_rx2_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx2_i(138)
  , pcs_m_comma_val              => cfg_rx2_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx2_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx2_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx2_i(115)
  , pcs_dec_bypass               => cfg_rx2_i(114)
  , pcs_el_buff_max_comp         => cfg_rx2_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx2_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx2_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx2_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx2_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx2_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx2_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx2_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx2_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx2_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx2_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx2_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx2_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx2_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx2_i(29)
  , pcs_buffers_bypass           => cfg_rx2_i(28)
  , pcs_sync_supported           => cfg_rx2_i(27)
  , pcs_replace_bypass           => cfg_rx2_i(26)
  , pcs_dscr_bypass              => cfg_rx2_i(25)
  , pcs_8b_dscr_sel              => cfg_rx2_i(24)
  , pcs_fsm_sel                  => cfg_rx2_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx2_i(21)
  , pma_pll_divm_en_n            => cfg_rx2_i(20)
  , pma_pll_divn_en_n            => cfg_rx2_i(19)
  , pma_cdr_cp                   => cfg_rx2_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx2_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx2_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx2_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx2_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx2_i(1)
  , pma_loopback                 => cfg_rx2_i(0)
  , location                     => location & ":CHANNEL3.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx2_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx2_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx2_ctrl_align_en_i
  , ALIGN_S_I => usr_rx2_ctrl_align_sync_i
  , REP_E_I   => usr_rx2_ctrl_replace_en_i
  , BUF_R_I   => usr_rx2_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx2_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx2_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx2_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx2_rst_n_i
  , CDR_R_I   => usr_rx2_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx2_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx2_pma_pll_rst_n_i

  , TST_I1    => usr_rx2_test_i(0)
  , TST_I2    => usr_rx2_test_i(1)
  , TST_I3    => usr_rx2_test_i(2)
  , TST_I4    => usr_rx2_test_i(3)

  , LOS_O     => usr_rx2_pma_loss_of_signal_o

  , DATA_O1   => usr_rx2_data_o(0)
  , DATA_O2   => usr_rx2_data_o(1)
  , DATA_O3   => usr_rx2_data_o(2)
  , DATA_O4   => usr_rx2_data_o(3)
  , DATA_O5   => usr_rx2_data_o(4)
  , DATA_O6   => usr_rx2_data_o(5)
  , DATA_O7   => usr_rx2_data_o(6)
  , DATA_O8   => usr_rx2_data_o(7)
  , DATA_O9   => usr_rx2_data_o(8)
  , DATA_O10  => usr_rx2_data_o(9)
  , DATA_O11  => usr_rx2_data_o(10)
  , DATA_O12  => usr_rx2_data_o(11)
  , DATA_O13  => usr_rx2_data_o(12)
  , DATA_O14  => usr_rx2_data_o(13)
  , DATA_O15  => usr_rx2_data_o(14)
  , DATA_O16  => usr_rx2_data_o(15)
  , DATA_O17  => usr_rx2_data_o(16)
  , DATA_O18  => usr_rx2_data_o(17)
  , DATA_O19  => usr_rx2_data_o(18)
  , DATA_O20  => usr_rx2_data_o(19)
  , DATA_O21  => usr_rx2_data_o(20)
  , DATA_O22  => usr_rx2_data_o(21)
  , DATA_O23  => usr_rx2_data_o(22)
  , DATA_O24  => usr_rx2_data_o(23)
  , DATA_O25  => usr_rx2_data_o(24)
  , DATA_O26  => usr_rx2_data_o(25)
  , DATA_O27  => usr_rx2_data_o(26)
  , DATA_O28  => usr_rx2_data_o(27)
  , DATA_O29  => usr_rx2_data_o(28)
  , DATA_O30  => usr_rx2_data_o(29)
  , DATA_O31  => usr_rx2_data_o(30)
  , DATA_O32  => usr_rx2_data_o(31)
  , DATA_O33  => usr_rx2_data_o(32)
  , DATA_O34  => usr_rx2_data_o(33)
  , DATA_O35  => usr_rx2_data_o(34)
  , DATA_O36  => usr_rx2_data_o(35)
  , DATA_O37  => usr_rx2_data_o(36)
  , DATA_O38  => usr_rx2_data_o(37)
  , DATA_O39  => usr_rx2_data_o(38)
  , DATA_O40  => usr_rx2_data_o(39)
  , DATA_O41  => usr_rx2_data_o(40)
  , DATA_O42  => usr_rx2_data_o(41)
  , DATA_O43  => usr_rx2_data_o(42)
  , DATA_O44  => usr_rx2_data_o(43)
  , DATA_O45  => usr_rx2_data_o(44)
  , DATA_O46  => usr_rx2_data_o(45)
  , DATA_O47  => usr_rx2_data_o(46)
  , DATA_O48  => usr_rx2_data_o(47)
  , DATA_O49  => usr_rx2_data_o(48)
  , DATA_O50  => usr_rx2_data_o(49)
  , DATA_O51  => usr_rx2_data_o(50)
  , DATA_O52  => usr_rx2_data_o(51)
  , DATA_O53  => usr_rx2_data_o(52)
  , DATA_O54  => usr_rx2_data_o(53)
  , DATA_O55  => usr_rx2_data_o(54)
  , DATA_O56  => usr_rx2_data_o(55)
  , DATA_O57  => usr_rx2_data_o(56)
  , DATA_O58  => usr_rx2_data_o(57)
  , DATA_O59  => usr_rx2_data_o(58)
  , DATA_O60  => usr_rx2_data_o(59)
  , DATA_O61  => usr_rx2_data_o(60)
  , DATA_O62  => usr_rx2_data_o(61)
  , DATA_O63  => usr_rx2_data_o(62)
  , DATA_O64  => usr_rx2_data_o(63)

  , CH_COM_O1 => usr_rx2_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx2_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx2_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx2_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx2_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx2_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx2_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx2_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx2_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx2_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx2_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx2_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx2_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx2_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx2_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx2_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx2_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx2_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx2_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx2_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx2_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx2_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx2_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx2_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx2_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx2_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx2_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx2_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx2_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx2_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx2_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx2_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx2_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx2_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx2_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx2_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx2_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx2_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx2_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx2_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx2_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx2_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx2_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx2_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx2_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx2_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx2_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx2_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx2_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx2_busy_o

  , TST_O1    => usr_rx2_test_o(0)
  , TST_O2    => usr_rx2_test_o(1)
  , TST_O3    => usr_rx2_test_o(2)
  , TST_O4    => usr_rx2_test_o(3)
  , TST_O5    => usr_rx2_test_o(4)
  , TST_O6    => usr_rx2_test_o(5)
  , TST_O7    => usr_rx2_test_o(6)
  , TST_O8    => usr_rx2_test_o(7)

  , LOCK_O    => usr_rx2_pll_lock_o

  , LINK      => LINK_RX2

  , RX_I      => pma_rx2_i
);
--#}}}#

-- txlane3: NX_CTX_L#{{{#
txlane3: NX_CTX_L generic map (
     pma_clk_pos          => cfg_tx3_i(31)
  ,  pcs_protocol_size    => cfg_tx3_i(30)
  ,  pcs_8b_scr_sel       => cfg_tx3_i(29)
  ,  pcs_scr_init         => cfg_tx3_i(28 downto 12)
  ,  pcs_scr_bypass       => cfg_tx3_i(11)
  ,  pcs_sync_supported   => cfg_tx3_i(10)
  ,  pcs_replace_bypass   => cfg_tx3_i(9)
  ,  pcs_enc_bypass       => cfg_tx3_i(8)
  ,  pcs_loopback         => cfg_tx3_i(7)
  ,  pcs_polarity         => cfg_tx3_i(6)
  ,  pcs_esistream_fsm_en => cfg_tx3_i(5)
  ,  test                 => cfg_tx3_i(4 downto 3)
  ,  pcs_bypass_pma_cdc   => cfg_tx3_i(2)
  ,  pcs_bypass_usr_cdc   => cfg_tx3_i(1)
  ,  pma_loopback         => cfg_tx3_i(0)
  ,  location             => location & ":CHANNEL4.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx3_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx3_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx3_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx3_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx3_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx3_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx3_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx3_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx3_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx3_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx3_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx3_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx3_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx3_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx3_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx3_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx3_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx3_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx3_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx3_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx3_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx3_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx3_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx3_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx3_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx3_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx3_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx3_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx3_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx3_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx3_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx3_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx3_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx3_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx3_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx3_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx3_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx3_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx3_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx3_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx3_ctrl_replace_en_i
  , RST_N_I  => usr_tx3_rst_n_i

  , TST_I1   => usr_tx3_test_i(0)
  , TST_I2   => usr_tx3_test_i(1)
  , TST_I3   => usr_tx3_test_i(2)
  , TST_I4   => usr_tx3_test_i(3)

  , DATA_I1  => usr_tx3_data_i(0)
  , DATA_I2  => usr_tx3_data_i(1)
  , DATA_I3  => usr_tx3_data_i(2)
  , DATA_I4  => usr_tx3_data_i(3)
  , DATA_I5  => usr_tx3_data_i(4)
  , DATA_I6  => usr_tx3_data_i(5)
  , DATA_I7  => usr_tx3_data_i(6)
  , DATA_I8  => usr_tx3_data_i(7)
  , DATA_I9  => usr_tx3_data_i(8)
  , DATA_I10 => usr_tx3_data_i(9)
  , DATA_I11 => usr_tx3_data_i(10)
  , DATA_I12 => usr_tx3_data_i(11)
  , DATA_I13 => usr_tx3_data_i(12)
  , DATA_I14 => usr_tx3_data_i(13)
  , DATA_I15 => usr_tx3_data_i(14)
  , DATA_I16 => usr_tx3_data_i(15)
  , DATA_I17 => usr_tx3_data_i(16)
  , DATA_I18 => usr_tx3_data_i(17)
  , DATA_I19 => usr_tx3_data_i(18)
  , DATA_I20 => usr_tx3_data_i(19)
  , DATA_I21 => usr_tx3_data_i(20)
  , DATA_I22 => usr_tx3_data_i(21)
  , DATA_I23 => usr_tx3_data_i(22)
  , DATA_I24 => usr_tx3_data_i(23)
  , DATA_I25 => usr_tx3_data_i(24)
  , DATA_I26 => usr_tx3_data_i(25)
  , DATA_I27 => usr_tx3_data_i(26)
  , DATA_I28 => usr_tx3_data_i(27)
  , DATA_I29 => usr_tx3_data_i(28)
  , DATA_I30 => usr_tx3_data_i(29)
  , DATA_I31 => usr_tx3_data_i(30)
  , DATA_I32 => usr_tx3_data_i(31)
  , DATA_I33 => usr_tx3_data_i(32)
  , DATA_I34 => usr_tx3_data_i(33)
  , DATA_I35 => usr_tx3_data_i(34)
  , DATA_I36 => usr_tx3_data_i(35)
  , DATA_I37 => usr_tx3_data_i(36)
  , DATA_I38 => usr_tx3_data_i(37)
  , DATA_I39 => usr_tx3_data_i(38)
  , DATA_I40 => usr_tx3_data_i(39)
  , DATA_I41 => usr_tx3_data_i(40)
  , DATA_I42 => usr_tx3_data_i(41)
  , DATA_I43 => usr_tx3_data_i(42)
  , DATA_I44 => usr_tx3_data_i(43)
  , DATA_I45 => usr_tx3_data_i(44)
  , DATA_I46 => usr_tx3_data_i(45)
  , DATA_I47 => usr_tx3_data_i(46)
  , DATA_I48 => usr_tx3_data_i(47)
  , DATA_I49 => usr_tx3_data_i(48)
  , DATA_I50 => usr_tx3_data_i(49)
  , DATA_I51 => usr_tx3_data_i(50)
  , DATA_I52 => usr_tx3_data_i(51)
  , DATA_I53 => usr_tx3_data_i(52)
  , DATA_I54 => usr_tx3_data_i(53)
  , DATA_I55 => usr_tx3_data_i(54)
  , DATA_I56 => usr_tx3_data_i(55)
  , DATA_I57 => usr_tx3_data_i(56)
  , DATA_I58 => usr_tx3_data_i(57)
  , DATA_I59 => usr_tx3_data_i(58)
  , DATA_I60 => usr_tx3_data_i(59)
  , DATA_I61 => usr_tx3_data_i(60)
  , DATA_I62 => usr_tx3_data_i(61)
  , DATA_I63 => usr_tx3_data_i(62)
  , DATA_I64 => usr_tx3_data_i(63)

  , TST_O1   => usr_tx3_test_o(0)
  , TST_O2   => usr_tx3_test_o(1)
  , TST_O3   => usr_tx3_test_o(2)
  , TST_O4   => usr_tx3_test_o(3)

  , BUSY_O   => usr_tx3_busy_o
  , CLK_E_I  => usr_tx3_pma_clk_en_i

  , LINK     => LINK_TX3

  , TX_O     => pma_tx3_o
);
--#}}}#

-- rxlane3: NX_CRX_L#{{{#
rxlane3: NX_CRX_L generic map (
    test                         => cfg_rx3_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx3_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx3_i(156)
  , pcs_debug_en                 => cfg_rx3_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx3_i(154)
  , pma_clk_pos                  => cfg_rx3_i(153)
  , pcs_protocol_size            => cfg_rx3_i(152)
  , pcs_loopback                 => cfg_rx3_i(151)
  , pcs_polarity                 => cfg_rx3_i(150)
  , pcs_p_comma_en               => cfg_rx3_i(149)
  , pcs_p_comma_val              => cfg_rx3_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx3_i(138)
  , pcs_m_comma_val              => cfg_rx3_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx3_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx3_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx3_i(115)
  , pcs_dec_bypass               => cfg_rx3_i(114)
  , pcs_el_buff_max_comp         => cfg_rx3_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx3_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx3_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx3_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx3_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx3_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx3_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx3_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx3_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx3_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx3_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx3_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx3_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx3_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx3_i(29)
  , pcs_buffers_bypass           => cfg_rx3_i(28)
  , pcs_sync_supported           => cfg_rx3_i(27)
  , pcs_replace_bypass           => cfg_rx3_i(26)
  , pcs_dscr_bypass              => cfg_rx3_i(25)
  , pcs_8b_dscr_sel              => cfg_rx3_i(24)
  , pcs_fsm_sel                  => cfg_rx3_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx3_i(21)
  , pma_pll_divm_en_n            => cfg_rx3_i(20)
  , pma_pll_divn_en_n            => cfg_rx3_i(19)
  , pma_cdr_cp                   => cfg_rx3_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx3_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx3_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx3_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx3_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx3_i(1)
  , pma_loopback                 => cfg_rx3_i(0)
  , location                     => location & ":CHANNEL4.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx3_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx3_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx3_ctrl_align_en_i
  , ALIGN_S_I => usr_rx3_ctrl_align_sync_i
  , REP_E_I   => usr_rx3_ctrl_replace_en_i
  , BUF_R_I   => usr_rx3_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx3_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx3_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx3_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx3_rst_n_i
  , CDR_R_I   => usr_rx3_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx3_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx3_pma_pll_rst_n_i

  , TST_I1    => usr_rx3_test_i(0)
  , TST_I2    => usr_rx3_test_i(1)
  , TST_I3    => usr_rx3_test_i(2)
  , TST_I4    => usr_rx3_test_i(3)

  , LOS_O     => usr_rx3_pma_loss_of_signal_o

  , DATA_O1   => usr_rx3_data_o(0)
  , DATA_O2   => usr_rx3_data_o(1)
  , DATA_O3   => usr_rx3_data_o(2)
  , DATA_O4   => usr_rx3_data_o(3)
  , DATA_O5   => usr_rx3_data_o(4)
  , DATA_O6   => usr_rx3_data_o(5)
  , DATA_O7   => usr_rx3_data_o(6)
  , DATA_O8   => usr_rx3_data_o(7)
  , DATA_O9   => usr_rx3_data_o(8)
  , DATA_O10  => usr_rx3_data_o(9)
  , DATA_O11  => usr_rx3_data_o(10)
  , DATA_O12  => usr_rx3_data_o(11)
  , DATA_O13  => usr_rx3_data_o(12)
  , DATA_O14  => usr_rx3_data_o(13)
  , DATA_O15  => usr_rx3_data_o(14)
  , DATA_O16  => usr_rx3_data_o(15)
  , DATA_O17  => usr_rx3_data_o(16)
  , DATA_O18  => usr_rx3_data_o(17)
  , DATA_O19  => usr_rx3_data_o(18)
  , DATA_O20  => usr_rx3_data_o(19)
  , DATA_O21  => usr_rx3_data_o(20)
  , DATA_O22  => usr_rx3_data_o(21)
  , DATA_O23  => usr_rx3_data_o(22)
  , DATA_O24  => usr_rx3_data_o(23)
  , DATA_O25  => usr_rx3_data_o(24)
  , DATA_O26  => usr_rx3_data_o(25)
  , DATA_O27  => usr_rx3_data_o(26)
  , DATA_O28  => usr_rx3_data_o(27)
  , DATA_O29  => usr_rx3_data_o(28)
  , DATA_O30  => usr_rx3_data_o(29)
  , DATA_O31  => usr_rx3_data_o(30)
  , DATA_O32  => usr_rx3_data_o(31)
  , DATA_O33  => usr_rx3_data_o(32)
  , DATA_O34  => usr_rx3_data_o(33)
  , DATA_O35  => usr_rx3_data_o(34)
  , DATA_O36  => usr_rx3_data_o(35)
  , DATA_O37  => usr_rx3_data_o(36)
  , DATA_O38  => usr_rx3_data_o(37)
  , DATA_O39  => usr_rx3_data_o(38)
  , DATA_O40  => usr_rx3_data_o(39)
  , DATA_O41  => usr_rx3_data_o(40)
  , DATA_O42  => usr_rx3_data_o(41)
  , DATA_O43  => usr_rx3_data_o(42)
  , DATA_O44  => usr_rx3_data_o(43)
  , DATA_O45  => usr_rx3_data_o(44)
  , DATA_O46  => usr_rx3_data_o(45)
  , DATA_O47  => usr_rx3_data_o(46)
  , DATA_O48  => usr_rx3_data_o(47)
  , DATA_O49  => usr_rx3_data_o(48)
  , DATA_O50  => usr_rx3_data_o(49)
  , DATA_O51  => usr_rx3_data_o(50)
  , DATA_O52  => usr_rx3_data_o(51)
  , DATA_O53  => usr_rx3_data_o(52)
  , DATA_O54  => usr_rx3_data_o(53)
  , DATA_O55  => usr_rx3_data_o(54)
  , DATA_O56  => usr_rx3_data_o(55)
  , DATA_O57  => usr_rx3_data_o(56)
  , DATA_O58  => usr_rx3_data_o(57)
  , DATA_O59  => usr_rx3_data_o(58)
  , DATA_O60  => usr_rx3_data_o(59)
  , DATA_O61  => usr_rx3_data_o(60)
  , DATA_O62  => usr_rx3_data_o(61)
  , DATA_O63  => usr_rx3_data_o(62)
  , DATA_O64  => usr_rx3_data_o(63)

  , CH_COM_O1 => usr_rx3_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx3_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx3_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx3_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx3_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx3_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx3_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx3_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx3_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx3_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx3_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx3_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx3_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx3_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx3_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx3_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx3_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx3_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx3_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx3_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx3_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx3_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx3_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx3_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx3_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx3_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx3_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx3_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx3_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx3_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx3_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx3_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx3_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx3_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx3_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx3_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx3_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx3_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx3_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx3_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx3_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx3_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx3_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx3_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx3_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx3_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx3_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx3_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx3_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx3_busy_o

  , TST_O1    => usr_rx3_test_o(0)
  , TST_O2    => usr_rx3_test_o(1)
  , TST_O3    => usr_rx3_test_o(2)
  , TST_O4    => usr_rx3_test_o(3)
  , TST_O5    => usr_rx3_test_o(4)
  , TST_O6    => usr_rx3_test_o(5)
  , TST_O7    => usr_rx3_test_o(6)
  , TST_O8    => usr_rx3_test_o(7)

  , LOCK_O    => usr_rx3_pll_lock_o

  , LINK      => LINK_RX3

  , RX_I      => pma_rx3_i
);
--#}}}#

-- txlane4: NX_CTX_L#{{{#
txlane4: NX_CTX_L generic map (
     pma_clk_pos          => cfg_tx4_i(31)
  ,  pcs_protocol_size    => cfg_tx4_i(30)
  ,  pcs_8b_scr_sel       => cfg_tx4_i(29)
  ,  pcs_scr_init         => cfg_tx4_i(28 downto 12)
  ,  pcs_scr_bypass       => cfg_tx4_i(11)
  ,  pcs_sync_supported   => cfg_tx4_i(10)
  ,  pcs_replace_bypass   => cfg_tx4_i(9)
  ,  pcs_enc_bypass       => cfg_tx4_i(8)
  ,  pcs_loopback         => cfg_tx4_i(7)
  ,  pcs_polarity         => cfg_tx4_i(6)
  ,  pcs_esistream_fsm_en => cfg_tx4_i(5)
  ,  test                 => cfg_tx4_i(4 downto 3)
  ,  pcs_bypass_pma_cdc   => cfg_tx4_i(2)
  ,  pcs_bypass_usr_cdc   => cfg_tx4_i(1)
  ,  pma_loopback         => cfg_tx4_i(0)
  ,  location             => location & ":CHANNEL5.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx4_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx4_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx4_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx4_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx4_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx4_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx4_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx4_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx4_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx4_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx4_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx4_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx4_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx4_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx4_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx4_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx4_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx4_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx4_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx4_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx4_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx4_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx4_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx4_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx4_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx4_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx4_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx4_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx4_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx4_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx4_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx4_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx4_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx4_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx4_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx4_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx4_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx4_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx4_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx4_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx4_ctrl_replace_en_i
  , RST_N_I  => usr_tx4_rst_n_i

  , TST_I1   => usr_tx4_test_i(0)
  , TST_I2   => usr_tx4_test_i(1)
  , TST_I3   => usr_tx4_test_i(2)
  , TST_I4   => usr_tx4_test_i(3)

  , DATA_I1  => usr_tx4_data_i(0)
  , DATA_I2  => usr_tx4_data_i(1)
  , DATA_I3  => usr_tx4_data_i(2)
  , DATA_I4  => usr_tx4_data_i(3)
  , DATA_I5  => usr_tx4_data_i(4)
  , DATA_I6  => usr_tx4_data_i(5)
  , DATA_I7  => usr_tx4_data_i(6)
  , DATA_I8  => usr_tx4_data_i(7)
  , DATA_I9  => usr_tx4_data_i(8)
  , DATA_I10 => usr_tx4_data_i(9)
  , DATA_I11 => usr_tx4_data_i(10)
  , DATA_I12 => usr_tx4_data_i(11)
  , DATA_I13 => usr_tx4_data_i(12)
  , DATA_I14 => usr_tx4_data_i(13)
  , DATA_I15 => usr_tx4_data_i(14)
  , DATA_I16 => usr_tx4_data_i(15)
  , DATA_I17 => usr_tx4_data_i(16)
  , DATA_I18 => usr_tx4_data_i(17)
  , DATA_I19 => usr_tx4_data_i(18)
  , DATA_I20 => usr_tx4_data_i(19)
  , DATA_I21 => usr_tx4_data_i(20)
  , DATA_I22 => usr_tx4_data_i(21)
  , DATA_I23 => usr_tx4_data_i(22)
  , DATA_I24 => usr_tx4_data_i(23)
  , DATA_I25 => usr_tx4_data_i(24)
  , DATA_I26 => usr_tx4_data_i(25)
  , DATA_I27 => usr_tx4_data_i(26)
  , DATA_I28 => usr_tx4_data_i(27)
  , DATA_I29 => usr_tx4_data_i(28)
  , DATA_I30 => usr_tx4_data_i(29)
  , DATA_I31 => usr_tx4_data_i(30)
  , DATA_I32 => usr_tx4_data_i(31)
  , DATA_I33 => usr_tx4_data_i(32)
  , DATA_I34 => usr_tx4_data_i(33)
  , DATA_I35 => usr_tx4_data_i(34)
  , DATA_I36 => usr_tx4_data_i(35)
  , DATA_I37 => usr_tx4_data_i(36)
  , DATA_I38 => usr_tx4_data_i(37)
  , DATA_I39 => usr_tx4_data_i(38)
  , DATA_I40 => usr_tx4_data_i(39)
  , DATA_I41 => usr_tx4_data_i(40)
  , DATA_I42 => usr_tx4_data_i(41)
  , DATA_I43 => usr_tx4_data_i(42)
  , DATA_I44 => usr_tx4_data_i(43)
  , DATA_I45 => usr_tx4_data_i(44)
  , DATA_I46 => usr_tx4_data_i(45)
  , DATA_I47 => usr_tx4_data_i(46)
  , DATA_I48 => usr_tx4_data_i(47)
  , DATA_I49 => usr_tx4_data_i(48)
  , DATA_I50 => usr_tx4_data_i(49)
  , DATA_I51 => usr_tx4_data_i(50)
  , DATA_I52 => usr_tx4_data_i(51)
  , DATA_I53 => usr_tx4_data_i(52)
  , DATA_I54 => usr_tx4_data_i(53)
  , DATA_I55 => usr_tx4_data_i(54)
  , DATA_I56 => usr_tx4_data_i(55)
  , DATA_I57 => usr_tx4_data_i(56)
  , DATA_I58 => usr_tx4_data_i(57)
  , DATA_I59 => usr_tx4_data_i(58)
  , DATA_I60 => usr_tx4_data_i(59)
  , DATA_I61 => usr_tx4_data_i(60)
  , DATA_I62 => usr_tx4_data_i(61)
  , DATA_I63 => usr_tx4_data_i(62)
  , DATA_I64 => usr_tx4_data_i(63)

  , TST_O1   => usr_tx4_test_o(0)
  , TST_O2   => usr_tx4_test_o(1)
  , TST_O3   => usr_tx4_test_o(2)
  , TST_O4   => usr_tx4_test_o(3)

  , BUSY_O   => usr_tx4_busy_o
  , CLK_E_I  => usr_tx4_pma_clk_en_i

  , LINK     => LINK_TX4

  , TX_O     => pma_tx4_o
);
--#}}}#

-- rxlane4: NX_CRX_L#{{{#
rxlane4: NX_CRX_L generic map (
    test                         => cfg_rx4_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx4_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx4_i(156)
  , pcs_debug_en                 => cfg_rx4_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx4_i(154)
  , pma_clk_pos                  => cfg_rx4_i(153)
  , pcs_protocol_size            => cfg_rx4_i(152)
  , pcs_loopback                 => cfg_rx4_i(151)
  , pcs_polarity                 => cfg_rx4_i(150)
  , pcs_p_comma_en               => cfg_rx4_i(149)
  , pcs_p_comma_val              => cfg_rx4_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx4_i(138)
  , pcs_m_comma_val              => cfg_rx4_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx4_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx4_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx4_i(115)
  , pcs_dec_bypass               => cfg_rx4_i(114)
  , pcs_el_buff_max_comp         => cfg_rx4_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx4_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx4_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx4_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx4_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx4_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx4_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx4_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx4_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx4_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx4_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx4_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx4_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx4_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx4_i(29)
  , pcs_buffers_bypass           => cfg_rx4_i(28)
  , pcs_sync_supported           => cfg_rx4_i(27)
  , pcs_replace_bypass           => cfg_rx4_i(26)
  , pcs_dscr_bypass              => cfg_rx4_i(25)
  , pcs_8b_dscr_sel              => cfg_rx4_i(24)
  , pcs_fsm_sel                  => cfg_rx4_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx4_i(21)
  , pma_pll_divm_en_n            => cfg_rx4_i(20)
  , pma_pll_divn_en_n            => cfg_rx4_i(19)
  , pma_cdr_cp                   => cfg_rx4_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx4_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx4_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx4_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx4_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx4_i(1)
  , pma_loopback                 => cfg_rx4_i(0)
  , location                     => location & ":CHANNEL5.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx4_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx4_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx4_ctrl_align_en_i
  , ALIGN_S_I => usr_rx4_ctrl_align_sync_i
  , REP_E_I   => usr_rx4_ctrl_replace_en_i
  , BUF_R_I   => usr_rx4_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx4_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx4_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx4_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx4_rst_n_i
  , CDR_R_I   => usr_rx4_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx4_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx4_pma_pll_rst_n_i

  , TST_I1    => usr_rx4_test_i(0)
  , TST_I2    => usr_rx4_test_i(1)
  , TST_I3    => usr_rx4_test_i(2)
  , TST_I4    => usr_rx4_test_i(3)

  , LOS_O     => usr_rx4_pma_loss_of_signal_o

  , DATA_O1   => usr_rx4_data_o(0)
  , DATA_O2   => usr_rx4_data_o(1)
  , DATA_O3   => usr_rx4_data_o(2)
  , DATA_O4   => usr_rx4_data_o(3)
  , DATA_O5   => usr_rx4_data_o(4)
  , DATA_O6   => usr_rx4_data_o(5)
  , DATA_O7   => usr_rx4_data_o(6)
  , DATA_O8   => usr_rx4_data_o(7)
  , DATA_O9   => usr_rx4_data_o(8)
  , DATA_O10  => usr_rx4_data_o(9)
  , DATA_O11  => usr_rx4_data_o(10)
  , DATA_O12  => usr_rx4_data_o(11)
  , DATA_O13  => usr_rx4_data_o(12)
  , DATA_O14  => usr_rx4_data_o(13)
  , DATA_O15  => usr_rx4_data_o(14)
  , DATA_O16  => usr_rx4_data_o(15)
  , DATA_O17  => usr_rx4_data_o(16)
  , DATA_O18  => usr_rx4_data_o(17)
  , DATA_O19  => usr_rx4_data_o(18)
  , DATA_O20  => usr_rx4_data_o(19)
  , DATA_O21  => usr_rx4_data_o(20)
  , DATA_O22  => usr_rx4_data_o(21)
  , DATA_O23  => usr_rx4_data_o(22)
  , DATA_O24  => usr_rx4_data_o(23)
  , DATA_O25  => usr_rx4_data_o(24)
  , DATA_O26  => usr_rx4_data_o(25)
  , DATA_O27  => usr_rx4_data_o(26)
  , DATA_O28  => usr_rx4_data_o(27)
  , DATA_O29  => usr_rx4_data_o(28)
  , DATA_O30  => usr_rx4_data_o(29)
  , DATA_O31  => usr_rx4_data_o(30)
  , DATA_O32  => usr_rx4_data_o(31)
  , DATA_O33  => usr_rx4_data_o(32)
  , DATA_O34  => usr_rx4_data_o(33)
  , DATA_O35  => usr_rx4_data_o(34)
  , DATA_O36  => usr_rx4_data_o(35)
  , DATA_O37  => usr_rx4_data_o(36)
  , DATA_O38  => usr_rx4_data_o(37)
  , DATA_O39  => usr_rx4_data_o(38)
  , DATA_O40  => usr_rx4_data_o(39)
  , DATA_O41  => usr_rx4_data_o(40)
  , DATA_O42  => usr_rx4_data_o(41)
  , DATA_O43  => usr_rx4_data_o(42)
  , DATA_O44  => usr_rx4_data_o(43)
  , DATA_O45  => usr_rx4_data_o(44)
  , DATA_O46  => usr_rx4_data_o(45)
  , DATA_O47  => usr_rx4_data_o(46)
  , DATA_O48  => usr_rx4_data_o(47)
  , DATA_O49  => usr_rx4_data_o(48)
  , DATA_O50  => usr_rx4_data_o(49)
  , DATA_O51  => usr_rx4_data_o(50)
  , DATA_O52  => usr_rx4_data_o(51)
  , DATA_O53  => usr_rx4_data_o(52)
  , DATA_O54  => usr_rx4_data_o(53)
  , DATA_O55  => usr_rx4_data_o(54)
  , DATA_O56  => usr_rx4_data_o(55)
  , DATA_O57  => usr_rx4_data_o(56)
  , DATA_O58  => usr_rx4_data_o(57)
  , DATA_O59  => usr_rx4_data_o(58)
  , DATA_O60  => usr_rx4_data_o(59)
  , DATA_O61  => usr_rx4_data_o(60)
  , DATA_O62  => usr_rx4_data_o(61)
  , DATA_O63  => usr_rx4_data_o(62)
  , DATA_O64  => usr_rx4_data_o(63)

  , CH_COM_O1 => usr_rx4_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx4_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx4_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx4_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx4_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx4_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx4_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx4_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx4_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx4_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx4_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx4_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx4_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx4_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx4_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx4_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx4_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx4_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx4_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx4_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx4_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx4_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx4_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx4_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx4_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx4_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx4_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx4_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx4_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx4_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx4_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx4_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx4_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx4_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx4_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx4_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx4_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx4_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx4_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx4_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx4_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx4_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx4_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx4_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx4_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx4_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx4_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx4_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx4_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx4_busy_o

  , TST_O1    => usr_rx4_test_o(0)
  , TST_O2    => usr_rx4_test_o(1)
  , TST_O3    => usr_rx4_test_o(2)
  , TST_O4    => usr_rx4_test_o(3)
  , TST_O5    => usr_rx4_test_o(4)
  , TST_O6    => usr_rx4_test_o(5)
  , TST_O7    => usr_rx4_test_o(6)
  , TST_O8    => usr_rx4_test_o(7)

  , LOCK_O    => usr_rx4_pll_lock_o

  , LINK      => LINK_RX4

  , RX_I      => pma_rx4_i
);
--#}}}#

-- txlane5: NX_CTX_L#{{{#
txlane5: NX_CTX_L generic map (
     pma_clk_pos          => cfg_tx5_i(31)
  ,  pcs_protocol_size    => cfg_tx5_i(30)
  ,  pcs_8b_scr_sel       => cfg_tx5_i(29)
  ,  pcs_scr_init         => cfg_tx5_i(28 downto 12)
  ,  pcs_scr_bypass       => cfg_tx5_i(11)
  ,  pcs_sync_supported   => cfg_tx5_i(10)
  ,  pcs_replace_bypass   => cfg_tx5_i(9)
  ,  pcs_enc_bypass       => cfg_tx5_i(8)
  ,  pcs_loopback         => cfg_tx5_i(7)
  ,  pcs_polarity         => cfg_tx5_i(6)
  ,  pcs_esistream_fsm_en => cfg_tx5_i(5)
  ,  test                 => cfg_tx5_i(4 downto 3)
  ,  pcs_bypass_pma_cdc   => cfg_tx5_i(2)
  ,  pcs_bypass_usr_cdc   => cfg_tx5_i(1)
  ,  pma_loopback         => cfg_tx5_i(0)
  ,  location             => location & ":CHANNEL6.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx5_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx5_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx5_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx5_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx5_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx5_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx5_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx5_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx5_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx5_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx5_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx5_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx5_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx5_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx5_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx5_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx5_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx5_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx5_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx5_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx5_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx5_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx5_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx5_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx5_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx5_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx5_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx5_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx5_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx5_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx5_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx5_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx5_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx5_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx5_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx5_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx5_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx5_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx5_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx5_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx5_ctrl_replace_en_i
  , RST_N_I  => usr_tx5_rst_n_i

  , TST_I1   => usr_tx5_test_i(0)
  , TST_I2   => usr_tx5_test_i(1)
  , TST_I3   => usr_tx5_test_i(2)
  , TST_I4   => usr_tx5_test_i(3)

  , DATA_I1  => usr_tx5_data_i(0)
  , DATA_I2  => usr_tx5_data_i(1)
  , DATA_I3  => usr_tx5_data_i(2)
  , DATA_I4  => usr_tx5_data_i(3)
  , DATA_I5  => usr_tx5_data_i(4)
  , DATA_I6  => usr_tx5_data_i(5)
  , DATA_I7  => usr_tx5_data_i(6)
  , DATA_I8  => usr_tx5_data_i(7)
  , DATA_I9  => usr_tx5_data_i(8)
  , DATA_I10 => usr_tx5_data_i(9)
  , DATA_I11 => usr_tx5_data_i(10)
  , DATA_I12 => usr_tx5_data_i(11)
  , DATA_I13 => usr_tx5_data_i(12)
  , DATA_I14 => usr_tx5_data_i(13)
  , DATA_I15 => usr_tx5_data_i(14)
  , DATA_I16 => usr_tx5_data_i(15)
  , DATA_I17 => usr_tx5_data_i(16)
  , DATA_I18 => usr_tx5_data_i(17)
  , DATA_I19 => usr_tx5_data_i(18)
  , DATA_I20 => usr_tx5_data_i(19)
  , DATA_I21 => usr_tx5_data_i(20)
  , DATA_I22 => usr_tx5_data_i(21)
  , DATA_I23 => usr_tx5_data_i(22)
  , DATA_I24 => usr_tx5_data_i(23)
  , DATA_I25 => usr_tx5_data_i(24)
  , DATA_I26 => usr_tx5_data_i(25)
  , DATA_I27 => usr_tx5_data_i(26)
  , DATA_I28 => usr_tx5_data_i(27)
  , DATA_I29 => usr_tx5_data_i(28)
  , DATA_I30 => usr_tx5_data_i(29)
  , DATA_I31 => usr_tx5_data_i(30)
  , DATA_I32 => usr_tx5_data_i(31)
  , DATA_I33 => usr_tx5_data_i(32)
  , DATA_I34 => usr_tx5_data_i(33)
  , DATA_I35 => usr_tx5_data_i(34)
  , DATA_I36 => usr_tx5_data_i(35)
  , DATA_I37 => usr_tx5_data_i(36)
  , DATA_I38 => usr_tx5_data_i(37)
  , DATA_I39 => usr_tx5_data_i(38)
  , DATA_I40 => usr_tx5_data_i(39)
  , DATA_I41 => usr_tx5_data_i(40)
  , DATA_I42 => usr_tx5_data_i(41)
  , DATA_I43 => usr_tx5_data_i(42)
  , DATA_I44 => usr_tx5_data_i(43)
  , DATA_I45 => usr_tx5_data_i(44)
  , DATA_I46 => usr_tx5_data_i(45)
  , DATA_I47 => usr_tx5_data_i(46)
  , DATA_I48 => usr_tx5_data_i(47)
  , DATA_I49 => usr_tx5_data_i(48)
  , DATA_I50 => usr_tx5_data_i(49)
  , DATA_I51 => usr_tx5_data_i(50)
  , DATA_I52 => usr_tx5_data_i(51)
  , DATA_I53 => usr_tx5_data_i(52)
  , DATA_I54 => usr_tx5_data_i(53)
  , DATA_I55 => usr_tx5_data_i(54)
  , DATA_I56 => usr_tx5_data_i(55)
  , DATA_I57 => usr_tx5_data_i(56)
  , DATA_I58 => usr_tx5_data_i(57)
  , DATA_I59 => usr_tx5_data_i(58)
  , DATA_I60 => usr_tx5_data_i(59)
  , DATA_I61 => usr_tx5_data_i(60)
  , DATA_I62 => usr_tx5_data_i(61)
  , DATA_I63 => usr_tx5_data_i(62)
  , DATA_I64 => usr_tx5_data_i(63)

  , TST_O1   => usr_tx5_test_o(0)
  , TST_O2   => usr_tx5_test_o(1)
  , TST_O3   => usr_tx5_test_o(2)
  , TST_O4   => usr_tx5_test_o(3)

  , BUSY_O   => usr_tx5_busy_o
  , CLK_E_I  => usr_tx5_pma_clk_en_i

  , LINK     => LINK_TX5

  , TX_O     => pma_tx5_o
);
--#}}}#

-- rxlane5: NX_CRX_L#{{{#
rxlane5: NX_CRX_L generic map (
    test                         => cfg_rx5_i(159 downto 158)
  , pcs_bypass_pma_cdc           => cfg_rx5_i(157)
  , pcs_bypass_usr_cdc           => cfg_rx5_i(156)
  , pcs_debug_en                 => cfg_rx5_i(155)
  , pcs_fsm_watchdog_en          => cfg_rx5_i(154)
  , pma_clk_pos                  => cfg_rx5_i(153)
  , pcs_protocol_size            => cfg_rx5_i(152)
  , pcs_loopback                 => cfg_rx5_i(151)
  , pcs_polarity                 => cfg_rx5_i(150)
  , pcs_p_comma_en               => cfg_rx5_i(149)
  , pcs_p_comma_val              => cfg_rx5_i(148 downto 139)
  , pcs_m_comma_en               => cfg_rx5_i(138)
  , pcs_m_comma_val              => cfg_rx5_i(137 downto 128)
  , pcs_comma_mask               => cfg_rx5_i(127 downto 118)
  , pcs_nb_comma_bef_realign     => cfg_rx5_i(117 downto 116)
  , pcs_align_bypass             => cfg_rx5_i(115)
  , pcs_dec_bypass               => cfg_rx5_i(114)
  , pcs_el_buff_max_comp         => cfg_rx5_i(113 downto 111)
  , pcs_el_buff_diff_bef_comp    => cfg_rx5_i(110 downto 108)
  , pcs_el_buff_only_one_skp     => cfg_rx5_i(107)
  , pcs_el_buff_underflow_handle => cfg_rx5_i(106)
  , pcs_el_buff_skp_seq_size     => cfg_rx5_i(105 downto 104)
  , pcs_el_buff_skp_char_0       => cfg_rx5_i(103 downto 95)
  , pcs_el_buff_skp_char_1       => cfg_rx5_i(94 downto 86)
  , pcs_el_buff_skp_char_2       => cfg_rx5_i(85 downto 77)
  , pcs_el_buff_skp_char_3       => cfg_rx5_i(76 downto 68)
  , pcs_el_buff_skp_header_size  => cfg_rx5_i(67 downto 66)
  , pcs_el_buff_skp_header_0     => cfg_rx5_i(65 downto 57)
  , pcs_el_buff_skp_header_1     => cfg_rx5_i(56 downto 48)
  , pcs_el_buff_skp_header_2     => cfg_rx5_i(47 downto 39)
  , pcs_el_buff_skp_header_3     => cfg_rx5_i(38 downto 30)
  , pcs_buffers_use_cdc          => cfg_rx5_i(29)
  , pcs_buffers_bypass           => cfg_rx5_i(28)
  , pcs_sync_supported           => cfg_rx5_i(27)
  , pcs_replace_bypass           => cfg_rx5_i(26)
  , pcs_dscr_bypass              => cfg_rx5_i(25)
  , pcs_8b_dscr_sel              => cfg_rx5_i(24)
  , pcs_fsm_sel                  => cfg_rx5_i(23 downto 22)
  , pma_pll_divf_en_n            => cfg_rx5_i(21)
  , pma_pll_divm_en_n            => cfg_rx5_i(20)
  , pma_pll_divn_en_n            => cfg_rx5_i(19)
  , pma_cdr_cp                   => cfg_rx5_i(18 downto 15)
  , pma_ctrl_term                => cfg_rx5_i(14 downto 9)
  , pma_pll_cpump_n              => cfg_rx5_i(8 downto 6)
  , pma_pll_divf                 => cfg_rx5_i(5 downto 4)
  , pma_pll_divm                 => cfg_rx5_i(3 downto 2)
  , pma_pll_divn                 => cfg_rx5_i(1)
  , pma_loopback                 => cfg_rx5_i(0)
  , location                     => location & ":CHANNEL6.CRX1"
 )
port map (
    DSCR_E_I  => usr_rx5_ctrl_dscr_en_i
  , DEC_E_I   => usr_rx5_ctrl_dec_en_i
  , ALIGN_E_I => usr_rx5_ctrl_align_en_i
  , ALIGN_S_I => usr_rx5_ctrl_align_sync_i
  , REP_E_I   => usr_rx5_ctrl_replace_en_i
  , BUF_R_I   => usr_rx5_ctrl_el_buff_rst_i

  , OVS_BS_I1 => usr_rx5_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2 => usr_rx5_ctrl_ovs_bit_sel_i(1)

  , BUF_FE_I  => usr_rx5_ctrl_el_buff_fifo_en_i
  , RST_N_I   => usr_rx5_rst_n_i
  , CDR_R_I   => usr_rx5_pma_cdr_rst_i
  , CKG_RN_I  => usr_rx5_pma_ckgen_rst_n_i
  , PLL_RN_I  => usr_rx5_pma_pll_rst_n_i

  , TST_I1    => usr_rx5_test_i(0)
  , TST_I2    => usr_rx5_test_i(1)
  , TST_I3    => usr_rx5_test_i(2)
  , TST_I4    => usr_rx5_test_i(3)

  , LOS_O     => usr_rx5_pma_loss_of_signal_o

  , DATA_O1   => usr_rx5_data_o(0)
  , DATA_O2   => usr_rx5_data_o(1)
  , DATA_O3   => usr_rx5_data_o(2)
  , DATA_O4   => usr_rx5_data_o(3)
  , DATA_O5   => usr_rx5_data_o(4)
  , DATA_O6   => usr_rx5_data_o(5)
  , DATA_O7   => usr_rx5_data_o(6)
  , DATA_O8   => usr_rx5_data_o(7)
  , DATA_O9   => usr_rx5_data_o(8)
  , DATA_O10  => usr_rx5_data_o(9)
  , DATA_O11  => usr_rx5_data_o(10)
  , DATA_O12  => usr_rx5_data_o(11)
  , DATA_O13  => usr_rx5_data_o(12)
  , DATA_O14  => usr_rx5_data_o(13)
  , DATA_O15  => usr_rx5_data_o(14)
  , DATA_O16  => usr_rx5_data_o(15)
  , DATA_O17  => usr_rx5_data_o(16)
  , DATA_O18  => usr_rx5_data_o(17)
  , DATA_O19  => usr_rx5_data_o(18)
  , DATA_O20  => usr_rx5_data_o(19)
  , DATA_O21  => usr_rx5_data_o(20)
  , DATA_O22  => usr_rx5_data_o(21)
  , DATA_O23  => usr_rx5_data_o(22)
  , DATA_O24  => usr_rx5_data_o(23)
  , DATA_O25  => usr_rx5_data_o(24)
  , DATA_O26  => usr_rx5_data_o(25)
  , DATA_O27  => usr_rx5_data_o(26)
  , DATA_O28  => usr_rx5_data_o(27)
  , DATA_O29  => usr_rx5_data_o(28)
  , DATA_O30  => usr_rx5_data_o(29)
  , DATA_O31  => usr_rx5_data_o(30)
  , DATA_O32  => usr_rx5_data_o(31)
  , DATA_O33  => usr_rx5_data_o(32)
  , DATA_O34  => usr_rx5_data_o(33)
  , DATA_O35  => usr_rx5_data_o(34)
  , DATA_O36  => usr_rx5_data_o(35)
  , DATA_O37  => usr_rx5_data_o(36)
  , DATA_O38  => usr_rx5_data_o(37)
  , DATA_O39  => usr_rx5_data_o(38)
  , DATA_O40  => usr_rx5_data_o(39)
  , DATA_O41  => usr_rx5_data_o(40)
  , DATA_O42  => usr_rx5_data_o(41)
  , DATA_O43  => usr_rx5_data_o(42)
  , DATA_O44  => usr_rx5_data_o(43)
  , DATA_O45  => usr_rx5_data_o(44)
  , DATA_O46  => usr_rx5_data_o(45)
  , DATA_O47  => usr_rx5_data_o(46)
  , DATA_O48  => usr_rx5_data_o(47)
  , DATA_O49  => usr_rx5_data_o(48)
  , DATA_O50  => usr_rx5_data_o(49)
  , DATA_O51  => usr_rx5_data_o(50)
  , DATA_O52  => usr_rx5_data_o(51)
  , DATA_O53  => usr_rx5_data_o(52)
  , DATA_O54  => usr_rx5_data_o(53)
  , DATA_O55  => usr_rx5_data_o(54)
  , DATA_O56  => usr_rx5_data_o(55)
  , DATA_O57  => usr_rx5_data_o(56)
  , DATA_O58  => usr_rx5_data_o(57)
  , DATA_O59  => usr_rx5_data_o(58)
  , DATA_O60  => usr_rx5_data_o(59)
  , DATA_O61  => usr_rx5_data_o(60)
  , DATA_O62  => usr_rx5_data_o(61)
  , DATA_O63  => usr_rx5_data_o(62)
  , DATA_O64  => usr_rx5_data_o(63)

  , CH_COM_O1 => usr_rx5_ctrl_char_is_comma_o(0)
  , CH_COM_O2 => usr_rx5_ctrl_char_is_comma_o(1)
  , CH_COM_O3 => usr_rx5_ctrl_char_is_comma_o(2)
  , CH_COM_O4 => usr_rx5_ctrl_char_is_comma_o(3)
  , CH_COM_O5 => usr_rx5_ctrl_char_is_comma_o(4)
  , CH_COM_O6 => usr_rx5_ctrl_char_is_comma_o(5)
  , CH_COM_O7 => usr_rx5_ctrl_char_is_comma_o(6)
  , CH_COM_O8 => usr_rx5_ctrl_char_is_comma_o(7)

  , CH_K_O1   => usr_rx5_ctrl_char_is_k_o(0)
  , CH_K_O2   => usr_rx5_ctrl_char_is_k_o(1)
  , CH_K_O3   => usr_rx5_ctrl_char_is_k_o(2)
  , CH_K_O4   => usr_rx5_ctrl_char_is_k_o(3)
  , CH_K_O5   => usr_rx5_ctrl_char_is_k_o(4)
  , CH_K_O6   => usr_rx5_ctrl_char_is_k_o(5)
  , CH_K_O7   => usr_rx5_ctrl_char_is_k_o(6)
  , CH_K_O8   => usr_rx5_ctrl_char_is_k_o(7)

  , NIT_O1    => usr_rx5_ctrl_not_in_table_o(0)
  , NIT_O2    => usr_rx5_ctrl_not_in_table_o(1)
  , NIT_O3    => usr_rx5_ctrl_not_in_table_o(2)
  , NIT_O4    => usr_rx5_ctrl_not_in_table_o(3)
  , NIT_O5    => usr_rx5_ctrl_not_in_table_o(4)
  , NIT_O6    => usr_rx5_ctrl_not_in_table_o(5)
  , NIT_O7    => usr_rx5_ctrl_not_in_table_o(6)
  , NIT_O8    => usr_rx5_ctrl_not_in_table_o(7)

  , D_ERR_O1  => usr_rx5_ctrl_disp_err_o(0)
  , D_ERR_O2  => usr_rx5_ctrl_disp_err_o(1)
  , D_ERR_O3  => usr_rx5_ctrl_disp_err_o(2)
  , D_ERR_O4  => usr_rx5_ctrl_disp_err_o(3)
  , D_ERR_O5  => usr_rx5_ctrl_disp_err_o(4)
  , D_ERR_O6  => usr_rx5_ctrl_disp_err_o(5)
  , D_ERR_O7  => usr_rx5_ctrl_disp_err_o(6)
  , D_ERR_O8  => usr_rx5_ctrl_disp_err_o(7)

  , CH_A_O1   => usr_rx5_ctrl_char_is_a_o(0)
  , CH_A_O2   => usr_rx5_ctrl_char_is_a_o(1)
  , CH_A_O3   => usr_rx5_ctrl_char_is_a_o(2)
  , CH_A_O4   => usr_rx5_ctrl_char_is_a_o(3)
  , CH_A_O5   => usr_rx5_ctrl_char_is_a_o(4)
  , CH_A_O6   => usr_rx5_ctrl_char_is_a_o(5)
  , CH_A_O7   => usr_rx5_ctrl_char_is_a_o(6)
  , CH_A_O8   => usr_rx5_ctrl_char_is_a_o(7)

  , CH_F_O1   => usr_rx5_ctrl_char_is_f_o(0)
  , CH_F_O2   => usr_rx5_ctrl_char_is_f_o(1)
  , CH_F_O3   => usr_rx5_ctrl_char_is_f_o(2)
  , CH_F_O4   => usr_rx5_ctrl_char_is_f_o(3)
  , CH_F_O5   => usr_rx5_ctrl_char_is_f_o(4)
  , CH_F_O6   => usr_rx5_ctrl_char_is_f_o(5)
  , CH_F_O7   => usr_rx5_ctrl_char_is_f_o(6)
  , CH_F_O8   => usr_rx5_ctrl_char_is_f_o(7)

  , ALIGN_O   => usr_rx5_ctrl_char_is_aligned_o
  , BUSY_O    => usr_rx5_busy_o

  , TST_O1    => usr_rx5_test_o(0)
  , TST_O2    => usr_rx5_test_o(1)
  , TST_O3    => usr_rx5_test_o(2)
  , TST_O4    => usr_rx5_test_o(3)
  , TST_O5    => usr_rx5_test_o(4)
  , TST_O6    => usr_rx5_test_o(5)
  , TST_O7    => usr_rx5_test_o(6)
  , TST_O8    => usr_rx5_test_o(7)

  , LOCK_O    => usr_rx5_pll_lock_o

  , LINK      => LINK_RX5

  , RX_I      => pma_rx5_i
);
--#}}}#

end NX_RTL;
--#}}}#
-- =================================================================================================
--   NX_PMA_L definition                                                                2018/11/30
-- =================================================================================================

-- NX_PMA_L#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_PMA_L is
 generic (
     main_test                   : bit_vector(7 downto 0) := (others => '0');
     rx_pma_half_step            : bit := '0';
     pll_pma_int_data_len        : bit := '0';
     pll_pma_cpump_n             : bit_vector(2 downto 0) := (others => '0');
     pll_pma_divf                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divm                : bit_vector(1 downto 0) := (others => '0');
     pll_pma_divn                : bit := '0';
     pll_pma_lvds_mux            : bit := '0';
     pll_pma_mux_ckref           : bit := '0';
     pll_pma_divf_en_n           : bit := '0';
     pll_pma_divm_en_n           : bit := '0';
     pll_pma_divn_en_n           : bit := '0';
     main_clk_to_fabric_div_mode : bit := '0';
     main_clk_to_fabric_div_en   : bit := '0';
     main_clk_to_fabric_sel      : bit := '0';
     main_use_only_usr_clock     : bit := '0';
     main_use_pcs_clk_2          : bit := '0';
     pcs_word_len                : bit_vector(1 downto 0) := (others => '0');
     pcs_ovs_mode                : bit := '0';
     pcs_pll_lock_count          : bit_vector(2 downto 0) := (others => '0');
     location                    : string := ""
 );
port (
    CLK_USER_I  : in  std_logic;
    CLK_REF_I   : in  std_logic;
--    CLK_I1      : in  std_logic;
--    CLK_I2      : in  std_logic;
--    CLK_I3      : in  std_logic;
--    CLK_I4      : in  std_logic;
--    CLK_I5      : in  std_logic;
--    CLK_I6      : in  std_logic;
--    CLK_I7      : in  std_logic;
--    CLK_I8      : in  std_logic;

    PRE_SG_I    : in  std_logic;
    PRE_EN_I    : in  std_logic;

    PRE_IS_I1   : in  std_logic;
    PRE_IS_I2   : in  std_logic;
    PRE_IS_I3   : in  std_logic;
    PRE_IS_I4   : in  std_logic;

    MAIN_SG_I   : in  std_logic;

    MAIN_EN_I1  : in  std_logic;
    MAIN_EN_I2  : in  std_logic;
    MAIN_EN_I3  : in  std_logic;
    MAIN_EN_I4  : in  std_logic;
    MAIN_EN_I5  : in  std_logic;
    MAIN_EN_I6  : in  std_logic;

    MARG_S_I1   : in  std_logic;
    MARG_S_I2   : in  std_logic;
    MARG_S_I3   : in  std_logic;
    MARG_S_I4   : in  std_logic;

    MARG_IS_I1  : in  std_logic;
    MARG_IS_I2  : in  std_logic;
    MARG_IS_I3  : in  std_logic;
    MARG_IS_I4  : in  std_logic;

    MARG_SV_I1  : in  std_logic;
    MARG_SV_I2  : in  std_logic;
    MARG_SV_I3  : in  std_logic;
    MARG_SV_I4  : in  std_logic;
    MARG_SV_I5  : in  std_logic;

    MARG_ISV_I1 : in  std_logic;
    MARG_ISV_I2 : in  std_logic;
    MARG_ISV_I3 : in  std_logic;
    MARG_ISV_I4 : in  std_logic;
    MARG_ISV_I5 : in  std_logic;

    POST_EN_I1  : in  std_logic;
    POST_EN_I2  : in  std_logic;
    POST_EN_I3  : in  std_logic;
    POST_EN_I4  : in  std_logic;
    POST_EN_I5  : in  std_logic;

    POST_SG_I   : in  std_logic;

    POST_IS_I1  : in  std_logic;
    POST_IS_I2  : in  std_logic;
    POST_IS_I3  : in  std_logic;
    POST_IS_I4  : in  std_logic;

    POST_ISV_I1 : in  std_logic;
    POST_ISV_I2 : in  std_logic;
    POST_ISV_I3 : in  std_logic;
    POST_ISV_I4 : in  std_logic;

    TX_SEL_I1   : in  std_logic;
    TX_SEL_I2   : in  std_logic;
    TX_SEL_I3   : in  std_logic;
    TX_SEL_I4   : in  std_logic;
    TX_SEL_I5   : in  std_logic;
    TX_SEL_I6   : in  std_logic;

    CT_CAP_I1   : in  std_logic;
    CT_CAP_I2   : in  std_logic;
    CT_CAP_I3   : in  std_logic;
    CT_CAP_I4   : in  std_logic;

    CT_RESP_I1  : in  std_logic;
    CT_RESP_I2  : in  std_logic;
    CT_RESP_I3  : in  std_logic;
    CT_RESP_I4  : in  std_logic;

    CT_RESN_I1  : in  std_logic;
    CT_RESN_I2  : in  std_logic;
    CT_RESN_I3  : in  std_logic;
    CT_RESN_I4  : in  std_logic;

    M_EYE_I     : in  std_logic;

    RX_SEL_I1   : in  std_logic;
    RX_SEL_I2   : in  std_logic;
    RX_SEL_I3   : in  std_logic;
    RX_SEL_I4   : in  std_logic;
    RX_SEL_I5   : in  std_logic;
    RX_SEL_I6   : in  std_logic;

    PLL_RN_I    : in  std_logic;
    RST_N_I     : in  std_logic;

    CAL_1P_I1   : in  std_logic;
    CAL_1P_I2   : in  std_logic;
    CAL_1P_I3   : in  std_logic;
    CAL_1P_I4   : in  std_logic;
    CAL_1P_I5   : in  std_logic;
    CAL_1P_I6   : in  std_logic;
    CAL_1P_I7   : in  std_logic;
    CAL_1P_I8   : in  std_logic;

    CAL_2N_I1   : in  std_logic;
    CAL_2N_I2   : in  std_logic;
    CAL_2N_I3   : in  std_logic;
    CAL_2N_I4   : in  std_logic;
    CAL_2N_I5   : in  std_logic;
    CAL_2N_I6   : in  std_logic;
    CAL_2N_I7   : in  std_logic;
    CAL_2N_I8   : in  std_logic;

    CAL_3N_I1   : in  std_logic;
    CAL_3N_I2   : in  std_logic;
    CAL_3N_I3   : in  std_logic;
    CAL_3N_I4   : in  std_logic;
    CAL_3N_I5   : in  std_logic;
    CAL_3N_I6   : in  std_logic;
    CAL_3N_I7   : in  std_logic;
    CAL_3N_I8   : in  std_logic;

    CAL_4P_I1   : in  std_logic;
    CAL_4P_I2   : in  std_logic;
    CAL_4P_I3   : in  std_logic;
    CAL_4P_I4   : in  std_logic;
    CAL_4P_I5   : in  std_logic;
    CAL_4P_I6   : in  std_logic;
    CAL_4P_I7   : in  std_logic;
    CAL_4P_I8   : in  std_logic;

    CAL_SEL_I1  : in  std_logic;
    CAL_SEL_I2  : in  std_logic;
    CAL_SEL_I3  : in  std_logic;
    CAL_SEL_I4  : in  std_logic;

    CAL_E_I     : in  std_logic;
    LOCK_E_I    : in  std_logic;
    OVS_E_I     : in  std_logic;

    TST_I1      : in  std_logic;
    TST_I2      : in  std_logic;
    TST_I3      : in  std_logic;
    TST_I4      : in  std_logic;
    TST_I5      : in  std_logic;
    TST_I6      : in  std_logic;
    TST_I7      : in  std_logic;
    TST_I8      : in  std_logic;

    CLK_O       : out std_logic;
    LOCK_O      : out std_logic;
    CAL_O       : out std_logic;

    TST_O1      : out std_logic;
    TST_O2      : out std_logic;
    TST_O3      : out std_logic;
    TST_O4      : out std_logic;
    TST_O5      : out std_logic;
    TST_O6      : out std_logic;
    TST_O7      : out std_logic;
    TST_O8      : out std_logic;

    LINK_TX0    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX1    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX2    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX3    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX4    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX5    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_RX0    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX1    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX2    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX3    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX4    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX5    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);

    CLK_EXT_I   : in  std_logic
);
end NX_PMA_L;
--#}}}#
-- =================================================================================================
--   NX_CRX_U definition                                                                2018/11/30
-- =================================================================================================

-- NX_CRX_U#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CRX_U is
 generic (
     cfg_rx_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_on_i                : bit := '0';
     cfg_rx_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_vref_sel_i                  : bit := '0';
     cfg_rx_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_divm_i                      : bit := '0';
     cfg_rx_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_loopback_i                      : bit := '0';
     cfg_rx_pma_clk_pos_i                       : bit := '0';
     cfg_rx_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divm_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divn_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divn_i                      : bit := '0';
     cfg_rx_pcs_debug_en_i                      : bit := '0';
     cfg_rx_pcs_bypass_pma_cdc_i                : bit := '0';
     cfg_rx_pcs_fsm_watchdog_en_i               : bit := '0';
     cfg_rx_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_polarity_i                      : bit := '0';
     cfg_rx_pcs_loopback_i                      : bit := '0';
     cfg_rx_pcs_dscr_bypass_i                   : bit := '0';
     cfg_rx_pcs_8b_dscr_sel_i                   : bit := '0';
     cfg_rx_pcs_replace_bypass_i                : bit := '0';
     cfg_rx_pcs_sync_supported_i                : bit := '0';
     cfg_rx_pcs_buffers_bypass_i                : bit := '0';
     cfg_rx_pcs_buffers_use_cdc_i               : bit := '0';
     cfg_rx_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_only_one_skp_i          : bit := '0';
     cfg_rx_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_dec_bypass_i                    : bit := '0';
     cfg_rx_pcs_align_bypass_i                  : bit := '0';
     cfg_rx_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_en_i                    : bit := '0';
     cfg_rx_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_p_comma_en_i                    : bit := '0';
     cfg_rx_pcs_bypass_usr_cdc_i                : bit := '0';
     cfg_rx_pcs_protocol_size_i                 : bit := '0';
     cfg_rx_gearbox_mode_i                      : bit := '0';
     cfg_rx_gearbox_en_i                        : bit := '0';
     location                     : string := ""
 );
port (
    DSCR_E_I  : in  std_logic;
    DEC_E_I   : in  std_logic;
    ALIGN_E_I : in  std_logic;
    ALIGN_S_I : in  std_logic;
    REP_E_I   : in  std_logic;
    BUF_R_I   : in  std_logic;

    OVS_BS_I1 : in  std_logic;
    OVS_BS_I2 : in  std_logic;

    RST_N_I   : in  std_logic;

    PMA_RSTN_I: in  std_logic;
    MEYE_RST_I: in  std_logic;
    PWDN_N_I  : in  std_logic;

    DBG_S_I1  : in  std_logic;
    DBG_S_I2  : in  std_logic;
    DBG_S_I3  : in  std_logic;

    DATA_O1   : out std_logic;
    DATA_O2   : out std_logic;
    DATA_O3   : out std_logic;
    DATA_O4   : out std_logic;
    DATA_O5   : out std_logic;
    DATA_O6   : out std_logic;
    DATA_O7   : out std_logic;
    DATA_O8   : out std_logic;
    DATA_O9   : out std_logic;
    DATA_O10  : out std_logic;
    DATA_O11  : out std_logic;
    DATA_O12  : out std_logic;
    DATA_O13  : out std_logic;
    DATA_O14  : out std_logic;
    DATA_O15  : out std_logic;
    DATA_O16  : out std_logic;
    DATA_O17  : out std_logic;
    DATA_O18  : out std_logic;
    DATA_O19  : out std_logic;
    DATA_O20  : out std_logic;
    DATA_O21  : out std_logic;
    DATA_O22  : out std_logic;
    DATA_O23  : out std_logic;
    DATA_O24  : out std_logic;
    DATA_O25  : out std_logic;
    DATA_O26  : out std_logic;
    DATA_O27  : out std_logic;
    DATA_O28  : out std_logic;
    DATA_O29  : out std_logic;
    DATA_O30  : out std_logic;
    DATA_O31  : out std_logic;
    DATA_O32  : out std_logic;
    DATA_O33  : out std_logic;
    DATA_O34  : out std_logic;
    DATA_O35  : out std_logic;
    DATA_O36  : out std_logic;
    DATA_O37  : out std_logic;
    DATA_O38  : out std_logic;
    DATA_O39  : out std_logic;
    DATA_O40  : out std_logic;
    DATA_O41  : out std_logic;
    DATA_O42  : out std_logic;
    DATA_O43  : out std_logic;
    DATA_O44  : out std_logic;
    DATA_O45  : out std_logic;
    DATA_O46  : out std_logic;
    DATA_O47  : out std_logic;
    DATA_O48  : out std_logic;
    DATA_O49  : out std_logic;
    DATA_O50  : out std_logic;
    DATA_O51  : out std_logic;
    DATA_O52  : out std_logic;
    DATA_O53  : out std_logic;
    DATA_O54  : out std_logic;
    DATA_O55  : out std_logic;
    DATA_O56  : out std_logic;
    DATA_O57  : out std_logic;
    DATA_O58  : out std_logic;
    DATA_O59  : out std_logic;
    DATA_O60  : out std_logic;
    DATA_O61  : out std_logic;
    DATA_O62  : out std_logic;
    DATA_O63  : out std_logic;
    DATA_O64  : out std_logic;

    CH_COM_O1 : out std_logic;
    CH_COM_O2 : out std_logic;
    CH_COM_O3 : out std_logic;
    CH_COM_O4 : out std_logic;
    CH_COM_O5 : out std_logic;
    CH_COM_O6 : out std_logic;
    CH_COM_O7 : out std_logic;
    CH_COM_O8 : out std_logic;

    CH_K_O1   : out std_logic;
    CH_K_O2   : out std_logic;
    CH_K_O3   : out std_logic;
    CH_K_O4   : out std_logic;
    CH_K_O5   : out std_logic;
    CH_K_O6   : out std_logic;
    CH_K_O7   : out std_logic;
    CH_K_O8   : out std_logic;

    NIT_O1    : out std_logic;
    NIT_O2    : out std_logic;
    NIT_O3    : out std_logic;
    NIT_O4    : out std_logic;
    NIT_O5    : out std_logic;
    NIT_O6    : out std_logic;
    NIT_O7    : out std_logic;
    NIT_O8    : out std_logic;

    D_ERR_O1  : out std_logic;
    D_ERR_O2  : out std_logic;
    D_ERR_O3  : out std_logic;
    D_ERR_O4  : out std_logic;
    D_ERR_O5  : out std_logic;
    D_ERR_O6  : out std_logic;
    D_ERR_O7  : out std_logic;
    D_ERR_O8  : out std_logic;

    CH_A_O1   : out std_logic;
    CH_A_O2   : out std_logic;
    CH_A_O3   : out std_logic;
    CH_A_O4   : out std_logic;
    CH_A_O5   : out std_logic;
    CH_A_O6   : out std_logic;
    CH_A_O7   : out std_logic;
    CH_A_O8   : out std_logic;

    CH_F_O1   : out std_logic;
    CH_F_O2   : out std_logic;
    CH_F_O3   : out std_logic;
    CH_F_O4   : out std_logic;
    CH_F_O5   : out std_logic;
    CH_F_O6   : out std_logic;
    CH_F_O7   : out std_logic;
    CH_F_O8   : out std_logic;

    ALIGN_O    : out std_logic;
    VREALIGN_O : out std_logic;
    BUSY_O     : out std_logic;

    TST_O1    : out std_logic;
    TST_O2    : out std_logic;
    TST_O3    : out std_logic;
    TST_O4    : out std_logic;
    TST_O5    : out std_logic;
    TST_O6    : out std_logic;
    TST_O7    : out std_logic;
    TST_O8    : out std_logic;

    LOS_O     : out std_logic;

    LL_FLOCK_O  : out std_logic;
    LL_SLOCK_O  : out std_logic;
    PLL_LOCK_O  : out std_logic;
    PLL_LOCKT_O : out std_logic;

    LINK      : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0)
);
end NX_CRX_U;
--#}}}#
-- =================================================================================================
--   NX_CTX_U definition                                                                2018/11/30
-- =================================================================================================

-- NX_CTX_U#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CTX_U is
 generic (
     cfg_tx_pcs_protocol_size_i    : bit := '0';
     cfg_tx_pcs_8b_scr_sel_i       : bit := '0';
     cfg_tx_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
     cfg_tx_pcs_scr_bypass_i       : bit := '0';
     cfg_tx_pcs_sync_supported_i   : bit := '0';
     cfg_tx_pcs_replace_bypass_i   : bit := '0';
     cfg_tx_pcs_enc_bypass_i       : bit := '0';
     cfg_tx_pcs_loopback_i         : bit := '0';
     cfg_tx_pcs_polarity_i         : bit := '0';
     cfg_tx_pcs_esistream_fsm_en_i : bit := '0';
     cfg_tx_pcs_bypass_pma_cdc_i   : bit := '0';
     cfg_tx_pcs_bypass_usr_cdc_i   : bit := '0';
     cfg_tx_pma_clk_pos_i          : bit := '0';
     cfg_tx_pma_loopback_i         : bit := '0';
     cfg_tx_gearbox_en_i           : bit := '0';
     cfg_tx_gearbox_mode_i         : bit := '0';

     location             : string := ""
 );
port (
    ENC_E_I1 : in  std_logic;
    ENC_E_I2 : in  std_logic;
    ENC_E_I3 : in  std_logic;
    ENC_E_I4 : in  std_logic;
    ENC_E_I5 : in  std_logic;
    ENC_E_I6 : in  std_logic;
    ENC_E_I7 : in  std_logic;
    ENC_E_I8 : in  std_logic;

    CH_K_I1  : in  std_logic;
    CH_K_I2  : in  std_logic;
    CH_K_I3  : in  std_logic;
    CH_K_I4  : in  std_logic;
    CH_K_I5  : in  std_logic;
    CH_K_I6  : in  std_logic;
    CH_K_I7  : in  std_logic;
    CH_K_I8  : in  std_logic;

    SCR_E_I1 : in  std_logic;
    SCR_E_I2 : in  std_logic;
    SCR_E_I3 : in  std_logic;
    SCR_E_I4 : in  std_logic;
    SCR_E_I5 : in  std_logic;
    SCR_E_I6 : in  std_logic;
    SCR_E_I7 : in  std_logic;
    SCR_E_I8 : in  std_logic;

    EOMF_I1  : in  std_logic;
    EOMF_I2  : in  std_logic;
    EOMF_I3  : in  std_logic;
    EOMF_I4  : in  std_logic;
    EOMF_I5  : in  std_logic;
    EOMF_I6  : in  std_logic;
    EOMF_I7  : in  std_logic;
    EOMF_I8  : in  std_logic;

    EOF_I1   : in  std_logic;
    EOF_I2   : in  std_logic;
    EOF_I3   : in  std_logic;
    EOF_I4   : in  std_logic;
    EOF_I5   : in  std_logic;
    EOF_I6   : in  std_logic;
    EOF_I7   : in  std_logic;
    EOF_I8   : in  std_logic;

    REP_E_I  : in  std_logic;
    RST_N_I  : in  std_logic;

    DATA_I1  : in  std_logic;
    DATA_I2  : in  std_logic;
    DATA_I3  : in  std_logic;
    DATA_I4  : in  std_logic;
    DATA_I5  : in  std_logic;
    DATA_I6  : in  std_logic;
    DATA_I7  : in  std_logic;
    DATA_I8  : in  std_logic;
    DATA_I9  : in  std_logic;
    DATA_I10 : in  std_logic;
    DATA_I11 : in  std_logic;
    DATA_I12 : in  std_logic;
    DATA_I13 : in  std_logic;
    DATA_I14 : in  std_logic;
    DATA_I15 : in  std_logic;
    DATA_I16 : in  std_logic;
    DATA_I17 : in  std_logic;
    DATA_I18 : in  std_logic;
    DATA_I19 : in  std_logic;
    DATA_I20 : in  std_logic;
    DATA_I21 : in  std_logic;
    DATA_I22 : in  std_logic;
    DATA_I23 : in  std_logic;
    DATA_I24 : in  std_logic;
    DATA_I25 : in  std_logic;
    DATA_I26 : in  std_logic;
    DATA_I27 : in  std_logic;
    DATA_I28 : in  std_logic;
    DATA_I29 : in  std_logic;
    DATA_I30 : in  std_logic;
    DATA_I31 : in  std_logic;
    DATA_I32 : in  std_logic;
    DATA_I33 : in  std_logic;
    DATA_I34 : in  std_logic;
    DATA_I35 : in  std_logic;
    DATA_I36 : in  std_logic;
    DATA_I37 : in  std_logic;
    DATA_I38 : in  std_logic;
    DATA_I39 : in  std_logic;
    DATA_I40 : in  std_logic;
    DATA_I41 : in  std_logic;
    DATA_I42 : in  std_logic;
    DATA_I43 : in  std_logic;
    DATA_I44 : in  std_logic;
    DATA_I45 : in  std_logic;
    DATA_I46 : in  std_logic;
    DATA_I47 : in  std_logic;
    DATA_I48 : in  std_logic;
    DATA_I49 : in  std_logic;
    DATA_I50 : in  std_logic;
    DATA_I51 : in  std_logic;
    DATA_I52 : in  std_logic;
    DATA_I53 : in  std_logic;
    DATA_I54 : in  std_logic;
    DATA_I55 : in  std_logic;
    DATA_I56 : in  std_logic;
    DATA_I57 : in  std_logic;
    DATA_I58 : in  std_logic;
    DATA_I59 : in  std_logic;
    DATA_I60 : in  std_logic;
    DATA_I61 : in  std_logic;
    DATA_I62 : in  std_logic;
    DATA_I63 : in  std_logic;
    DATA_I64 : in  std_logic;

    BUSY_O   : out std_logic;
    INV_K_O  : out std_logic;

    PWDN_N_I : in  std_logic;
    CLK_E_I  : in  std_logic;

    CLK_O    : out std_logic;

    LINK     : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0)
);
end NX_CTX_U;
--#}}}#
-- =================================================================================================
--   NX_HSSL_U_FULL declaration                                                          2019/06/20
-- =================================================================================================

-- NX_HSSL_U_FULL#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_HSSL_U_FULL is
generic (
   -- PMA
   cfg_pll_pma_int_data_len_i            : bit := '0';
   cfg_pll_pma_cpump_i                   : bit_vector( 3 downto 0) := (others => '0');
   cfg_pll_pma_divl_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_divm_i                    : bit := '0';
   cfg_pll_pma_divn_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_lvds_en_i                 : bit := '0';
   cfg_pll_pma_lvds_mux_i                : bit := '0';
   cfg_pll_pma_mux_ckref_i               : bit := '0';
   cfg_pll_pma_gbx_en_i                  : bit := '0';
   cfg_pll_pma_ckref_ext_i               : bit := '0';
   cfg_main_clk_to_fabric_div_mode_i     : bit := '0';
   cfg_main_clk_to_fabric_div_en_i       : bit := '0';
   cfg_main_clk_to_fabric_sel_i          : bit := '0';
   cfg_main_rclk_to_fabric_sel_i         : bit_vector( 1 downto 0) := (others => '0');
   cfg_main_use_only_usr_clock_i         : bit := '0';
   tx_usrclk_use_pcs_clk_2               : bit := '0';
   rx_usrclk_use_pcs_clk_2               : bit := '0';
   cfg_pcs_word_len_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pcs_ovs_en_i                      : bit := '0';
   cfg_pcs_ovs_mode_i                    : bit := '0';
   cfg_pcs_pll_lock_ppm_i                : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_m_eye_i            : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_up_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_dn_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_coarse_ena_i : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_fine_ena_i   : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_step_i       : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_mode_i        : bit_vector( 1 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_locked_i      : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_unlocked_i    : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_1        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_2        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx1_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx2_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx3_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx0_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx1_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx2_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx3_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx0_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_test_mode_i                       : bit_vector( 1 downto 0) := (others => '0');

   --LANE 0
   --TX
   cfg_tx0_pcs_protocol_size_i    : bit := '0';
   cfg_tx0_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx0_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx0_pcs_scr_bypass_i       : bit := '0';
   cfg_tx0_pcs_sync_supported_i   : bit := '0';
   cfg_tx0_pcs_replace_bypass_i   : bit := '0';
   cfg_tx0_pcs_enc_bypass_i       : bit := '0';
   cfg_tx0_pcs_loopback_i         : bit := '0';
   cfg_tx0_pcs_polarity_i         : bit := '0';
   cfg_tx0_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx0_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx0_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx0_pma_clk_pos_i          : bit := '0';
   cfg_tx0_pma_loopback_i         : bit := '0';
   cfg_tx0_gearbox_en_i           : bit := '0';
   cfg_tx0_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx0_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_peak_detect_on_i                : bit := '0';
   cfg_rx0_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx0_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_dco_divm_i                      : bit := '0';
   cfg_rx0_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_loopback_i                      : bit := '0';
   cfg_rx0_pma_clk_pos_i                       : bit := '0';
   cfg_rx0_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx0_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pma_pll_divn_i                      : bit := '0';
   cfg_rx0_pcs_debug_en_i                      : bit := '0';
   cfg_rx0_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx0_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx0_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_polarity_i                      : bit := '0';
   cfg_rx0_pcs_loopback_i                      : bit := '0';
   cfg_rx0_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx0_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx0_pcs_replace_bypass_i                : bit := '0';
   cfg_rx0_pcs_sync_supported_i                : bit := '0';
   cfg_rx0_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx0_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx0_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx0_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx0_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx0_pcs_align_bypass_i                  : bit := '0';
   cfg_rx0_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx0_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx0_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx0_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx0_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx0_pcs_protocol_size_i                 : bit := '0';
   cfg_rx0_gearbox_mode_i                      : bit := '0';
   cfg_rx0_gearbox_en_i                        : bit := '0';

   --LANE 1
   --TX
   cfg_tx1_pcs_protocol_size_i    : bit := '0';
   cfg_tx1_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx1_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx1_pcs_scr_bypass_i       : bit := '0';
   cfg_tx1_pcs_sync_supported_i   : bit := '0';
   cfg_tx1_pcs_replace_bypass_i   : bit := '0';
   cfg_tx1_pcs_enc_bypass_i       : bit := '0';
   cfg_tx1_pcs_loopback_i         : bit := '0';
   cfg_tx1_pcs_polarity_i         : bit := '0';
   cfg_tx1_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx1_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx1_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx1_pma_clk_pos_i          : bit := '0';
   cfg_tx1_pma_loopback_i         : bit := '0';
   cfg_tx1_gearbox_en_i           : bit := '0';
   cfg_tx1_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx1_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_peak_detect_on_i                : bit := '0';
   cfg_rx1_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx1_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_dco_divm_i                      : bit := '0';
   cfg_rx1_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_loopback_i                      : bit := '0';
   cfg_rx1_pma_clk_pos_i                       : bit := '0';
   cfg_rx1_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx1_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pma_pll_divn_i                      : bit := '0';
   cfg_rx1_pcs_debug_en_i                      : bit := '0';
   cfg_rx1_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx1_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx1_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_polarity_i                      : bit := '0';
   cfg_rx1_pcs_loopback_i                      : bit := '0';
   cfg_rx1_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx1_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx1_pcs_replace_bypass_i                : bit := '0';
   cfg_rx1_pcs_sync_supported_i                : bit := '0';
   cfg_rx1_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx1_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx1_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx1_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx1_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx1_pcs_align_bypass_i                  : bit := '0';
   cfg_rx1_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx1_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx1_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx1_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx1_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx1_pcs_protocol_size_i                 : bit := '0';
   cfg_rx1_gearbox_mode_i                      : bit := '0';
   cfg_rx1_gearbox_en_i                        : bit := '0';

   --LANE 2
   --TX
   cfg_tx2_pcs_protocol_size_i    : bit := '0';
   cfg_tx2_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx2_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx2_pcs_scr_bypass_i       : bit := '0';
   cfg_tx2_pcs_sync_supported_i   : bit := '0';
   cfg_tx2_pcs_replace_bypass_i   : bit := '0';
   cfg_tx2_pcs_enc_bypass_i       : bit := '0';
   cfg_tx2_pcs_loopback_i         : bit := '0';
   cfg_tx2_pcs_polarity_i         : bit := '0';
   cfg_tx2_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx2_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx2_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx2_pma_clk_pos_i          : bit := '0';
   cfg_tx2_pma_loopback_i         : bit := '0';
   cfg_tx2_gearbox_en_i           : bit := '0';
   cfg_tx2_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx2_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_peak_detect_on_i                : bit := '0';
   cfg_rx2_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx2_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_dco_divm_i                      : bit := '0';
   cfg_rx2_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_loopback_i                      : bit := '0';
   cfg_rx2_pma_clk_pos_i                       : bit := '0';
   cfg_rx2_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx2_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pma_pll_divn_i                      : bit := '0';
   cfg_rx2_pcs_debug_en_i                      : bit := '0';
   cfg_rx2_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx2_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx2_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_polarity_i                      : bit := '0';
   cfg_rx2_pcs_loopback_i                      : bit := '0';
   cfg_rx2_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx2_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx2_pcs_replace_bypass_i                : bit := '0';
   cfg_rx2_pcs_sync_supported_i                : bit := '0';
   cfg_rx2_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx2_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx2_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx2_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx2_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx2_pcs_align_bypass_i                  : bit := '0';
   cfg_rx2_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx2_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx2_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx2_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx2_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx2_pcs_protocol_size_i                 : bit := '0';
   cfg_rx2_gearbox_mode_i                      : bit := '0';
   cfg_rx2_gearbox_en_i                        : bit := '0';

   --LANE 3
   --TX
   cfg_tx3_pcs_protocol_size_i    : bit := '0';
   cfg_tx3_pcs_8b_scr_sel_i       : bit := '0';
   cfg_tx3_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
   cfg_tx3_pcs_scr_bypass_i       : bit := '0';
   cfg_tx3_pcs_sync_supported_i   : bit := '0';
   cfg_tx3_pcs_replace_bypass_i   : bit := '0';
   cfg_tx3_pcs_enc_bypass_i       : bit := '0';
   cfg_tx3_pcs_loopback_i         : bit := '0';
   cfg_tx3_pcs_polarity_i         : bit := '0';
   cfg_tx3_pcs_esistream_fsm_en_i : bit := '0';
   cfg_tx3_pcs_bypass_pma_cdc_i   : bit := '0';
   cfg_tx3_pcs_bypass_usr_cdc_i   : bit := '0';
   cfg_tx3_pma_clk_pos_i          : bit := '0';
   cfg_tx3_pma_loopback_i         : bit := '0';
   cfg_tx3_gearbox_en_i           : bit := '0';
   cfg_tx3_gearbox_mode_i         : bit := '0';
   --RX
   cfg_rx3_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_peak_detect_on_i                : bit := '0';
   cfg_rx3_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_dco_vref_sel_i                  : bit := '0';
   cfg_rx3_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_dco_divm_i                      : bit := '0';
   cfg_rx3_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_loopback_i                      : bit := '0';
   cfg_rx3_pma_clk_pos_i                       : bit := '0';
   cfg_rx3_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divf_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_divm_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_divn_en_n_i                 : bit := '0';
   cfg_rx3_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pma_pll_divn_i                      : bit := '0';
   cfg_rx3_pcs_debug_en_i                      : bit := '0';
   cfg_rx3_pcs_bypass_pma_cdc_i                : bit := '0';
   cfg_rx3_pcs_fsm_watchdog_en_i               : bit := '0';
   cfg_rx3_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_polarity_i                      : bit := '0';
   cfg_rx3_pcs_loopback_i                      : bit := '0';
   cfg_rx3_pcs_dscr_bypass_i                   : bit := '0';
   cfg_rx3_pcs_8b_dscr_sel_i                   : bit := '0';
   cfg_rx3_pcs_replace_bypass_i                : bit := '0';
   cfg_rx3_pcs_sync_supported_i                : bit := '0';
   cfg_rx3_pcs_buffers_bypass_i                : bit := '0';
   cfg_rx3_pcs_buffers_use_cdc_i               : bit := '0';
   cfg_rx3_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_only_one_skp_i          : bit := '0';
   cfg_rx3_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
   cfg_rx3_pcs_dec_bypass_i                    : bit := '0';
   cfg_rx3_pcs_align_bypass_i                  : bit := '0';
   cfg_rx3_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
   cfg_rx3_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_m_comma_en_i                    : bit := '0';
   cfg_rx3_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
   cfg_rx3_pcs_p_comma_en_i                    : bit := '0';
   cfg_rx3_pcs_bypass_usr_cdc_i                : bit := '0';
   cfg_rx3_pcs_protocol_size_i                 : bit := '0';
   cfg_rx3_gearbox_mode_i                      : bit := '0';
   cfg_rx3_gearbox_en_i                        : bit := '0';

   location   : string := ""
 );
port (
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ MAIN ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- PMA
   hssl_clk_user_tx_i                     : in  std_logic;
   hssl_clk_user_rx_i                     : in  std_logic;
   hssl_clk_ref_i                         : in  std_logic;
   hssl_clock_o                           : out std_logic;
   hssl_rclock_o                          : out std_logic;
   usr_dyn_cfg_en_i                       : in  std_logic;
   usr_dyn_cfg_lane_cs_n_i                : in  std_logic_vector(3 downto 0);
   usr_dyn_cfg_calibration_cs_n_i         : in  std_logic;
   usr_dyn_cfg_we_n_i                     : in  std_logic;
   usr_dyn_cfg_addr_i                     : in  std_logic_vector(3 downto 0);
   usr_dyn_cfg_wdata_sel_i                : in  std_logic;
   usr_dyn_cfg_wdata_i                    : in  std_logic_vector(11 downto 0);
   usr_pll_pma_rst_n_i                    : in  std_logic;
   usr_pll_pma_pwr_down_n_i               : in  std_logic;
   usr_main_rst_n_i                       : in  std_logic;
   usr_pll_lock_o                         : out std_logic;
   usr_pll_pma_lock_analog_o              : out std_logic;
   usr_pll_ckfb_lock_o                    : out std_logic;
   usr_calibrate_pma_out_o                : out std_logic;
   usr_main_async_debug_lane_sel_i        : in  std_logic_vector(1 downto 0);
   usr_main_async_debug_ack_i             : in  std_logic;
   usr_main_async_debug_req_o             : out std_logic;
   usr_main_rx_pma_ll_out_o               : out std_logic_vector(19 downto 0);
   scan_en_i                              : in  std_logic;
   scan_in_i                              : in  std_logic_vector(7 downto 0);
   scan_out_o                             : out std_logic_vector(7 downto 0);


   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 0 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
   usr_tx0_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx0_ctrl_replace_en_i        : in  std_logic;
   usr_tx0_rst_n_i                  : in  std_logic;
   usr_tx0_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx0_busy_o                   : out std_logic;
   usr_tx0_ctrl_invalid_k_o         : out std_logic;
   usr_tx0_ctrl_driver_pwrdwn_n_i   : in  std_logic;
   usr_tx0_pma_clk_en_i             : in  std_logic;
   usr_tx0_pma_tx_clk_o             : out std_logic;

    -- RX - Fabric Interface
   usr_rx0_ctrl_dscr_en_i         : in  std_logic;
   usr_rx0_ctrl_dec_en_i          : in  std_logic;
   usr_rx0_ctrl_align_en_i        : in  std_logic;
   usr_rx0_ctrl_align_sync_i      : in  std_logic;
   usr_rx0_ctrl_replace_en_i      : in  std_logic;
   usr_rx0_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx0_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx0_rst_n_i                : in  std_logic;
   usr_rx0_pma_rst_n_i            : in  std_logic;
   usr_rx0_pma_m_eye_rst_i        : in  std_logic;
   usr_rx0_pma_pwr_down_n_i       : in  std_logic;
   usr_rx0_ctrl_debug_sel_i       : in  std_logic_vector(2 downto 0);
   usr_rx0_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx0_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx0_ctrl_char_is_aligned_o : out std_logic;
   usr_rx0_ctrl_valid_realign_o   : out std_logic;
   usr_rx0_busy_o                 : out std_logic;
   usr_rx0_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx0_pma_loss_of_signal_o   : out std_logic;
   usr_rx0_pma_ll_fast_locked_o   : out std_logic;
   usr_rx0_pma_ll_slow_locked_o   : out std_logic;
   usr_rx0_pma_pll_lock_o         : out std_logic;
   usr_rx0_pma_pll_lock_track_o   : out std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 1 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
   usr_tx1_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx1_ctrl_replace_en_i        : in  std_logic;
   usr_tx1_rst_n_i                  : in  std_logic;
   usr_tx1_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx1_busy_o                   : out std_logic;
   usr_tx1_ctrl_invalid_k_o         : out std_logic;
   usr_tx1_ctrl_driver_pwrdwn_n_i   : in  std_logic;
   usr_tx1_pma_clk_en_i             : in  std_logic;
   usr_tx1_pma_tx_clk_o             : out std_logic;

    -- RX - Fabric Interface
   usr_rx1_ctrl_dscr_en_i         : in  std_logic;
   usr_rx1_ctrl_dec_en_i          : in  std_logic;
   usr_rx1_ctrl_align_en_i        : in  std_logic;
   usr_rx1_ctrl_align_sync_i      : in  std_logic;
   usr_rx1_ctrl_replace_en_i      : in  std_logic;
   usr_rx1_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx1_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx1_rst_n_i                : in  std_logic;
   usr_rx1_pma_rst_n_i            : in  std_logic;
   usr_rx1_pma_m_eye_rst_i        : in  std_logic;
   usr_rx1_pma_pwr_down_n_i       : in  std_logic;
   usr_rx1_ctrl_debug_sel_i       : in  std_logic_vector(2 downto 0);
   usr_rx1_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx1_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx1_ctrl_char_is_aligned_o : out std_logic;
   usr_rx1_ctrl_valid_realign_o   : out std_logic;
   usr_rx1_busy_o                 : out std_logic;
   usr_rx1_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx1_pma_loss_of_signal_o   : out std_logic;
   usr_rx1_pma_ll_fast_locked_o   : out std_logic;
   usr_rx1_pma_ll_slow_locked_o   : out std_logic;
   usr_rx1_pma_pll_lock_o         : out std_logic;
   usr_rx1_pma_pll_lock_track_o   : out std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 2 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
   usr_tx2_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx2_ctrl_replace_en_i        : in  std_logic;
   usr_tx2_rst_n_i                  : in  std_logic;
   usr_tx2_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx2_busy_o                   : out std_logic;
   usr_tx2_ctrl_invalid_k_o         : out std_logic;
   usr_tx2_ctrl_driver_pwrdwn_n_i   : in  std_logic;
   usr_tx2_pma_clk_en_i             : in  std_logic;
   usr_tx2_pma_tx_clk_o             : out std_logic;

   -- RX - Fabric Interface
   usr_rx2_ctrl_dscr_en_i         : in  std_logic;
   usr_rx2_ctrl_dec_en_i          : in  std_logic;
   usr_rx2_ctrl_align_en_i        : in  std_logic;
   usr_rx2_ctrl_align_sync_i      : in  std_logic;
   usr_rx2_ctrl_replace_en_i      : in  std_logic;
   usr_rx2_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx2_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx2_rst_n_i                : in  std_logic;
   usr_rx2_pma_rst_n_i            : in  std_logic;
   usr_rx2_pma_m_eye_rst_i        : in  std_logic;
   usr_rx2_pma_pwr_down_n_i       : in  std_logic;
   usr_rx2_ctrl_debug_sel_i       : in  std_logic_vector(2 downto 0);
   usr_rx2_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx2_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx2_ctrl_char_is_aligned_o : out std_logic;
   usr_rx2_ctrl_valid_realign_o   : out std_logic;
   usr_rx2_busy_o                 : out std_logic;
   usr_rx2_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx2_pma_loss_of_signal_o   : out std_logic;
   usr_rx2_pma_ll_fast_locked_o   : out std_logic;
   usr_rx2_pma_ll_slow_locked_o   : out std_logic;
   usr_rx2_pma_pll_lock_o         : out std_logic;
   usr_rx2_pma_pll_lock_track_o   : out std_logic;

   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   --~~~ LANE 3 ~~~
   --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
   -- TX - Fabric Interface
   usr_tx3_ctrl_enc_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_char_is_k_i         : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_scr_en_i            : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_end_of_multiframe_i : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_end_of_frame_i      : in  std_logic_vector(7 downto 0);
   usr_tx3_ctrl_replace_en_i        : in  std_logic;
   usr_tx3_rst_n_i                  : in  std_logic;
   usr_tx3_data_i                   : in  std_logic_vector(63 downto 0);
   usr_tx3_busy_o                   : out std_logic;
   usr_tx3_ctrl_invalid_k_o         : out std_logic;
   usr_tx3_ctrl_driver_pwrdwn_n_i   : in  std_logic;
   usr_tx3_pma_clk_en_i             : in  std_logic;
   usr_tx3_pma_tx_clk_o             : out std_logic;

   -- RX - Fabric Interface
   usr_rx3_ctrl_dscr_en_i         : in  std_logic;
   usr_rx3_ctrl_dec_en_i          : in  std_logic;
   usr_rx3_ctrl_align_en_i        : in  std_logic;
   usr_rx3_ctrl_align_sync_i      : in  std_logic;
   usr_rx3_ctrl_replace_en_i      : in  std_logic;
   usr_rx3_ctrl_el_buff_rst_i     : in  std_logic;
   usr_rx3_ctrl_ovs_bit_sel_i     : in  std_logic_vector(1 downto 0);
   usr_rx3_rst_n_i                : in  std_logic;
   usr_rx3_pma_rst_n_i            : in  std_logic;
   usr_rx3_pma_m_eye_rst_i        : in  std_logic;
   usr_rx3_pma_pwr_down_n_i       : in  std_logic;
   usr_rx3_ctrl_debug_sel_i       : in  std_logic_vector(2 downto 0);
   usr_rx3_data_o                 : out std_logic_vector(63 downto 0);
   usr_rx3_ctrl_char_is_comma_o   : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_k_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_not_in_table_o    : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_disp_err_o        : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_a_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_f_o       : out std_logic_vector(7 downto 0);
   usr_rx3_ctrl_char_is_aligned_o : out std_logic;
   usr_rx3_ctrl_valid_realign_o   : out std_logic;
   usr_rx3_busy_o                 : out std_logic;
   usr_rx3_test_o                 : out std_logic_vector(7 downto 0);
   usr_rx3_pma_loss_of_signal_o   : out std_logic;
   usr_rx3_pma_ll_fast_locked_o   : out std_logic;
   usr_rx3_pma_ll_slow_locked_o   : out std_logic;
   usr_rx3_pma_pll_lock_o         : out std_logic;
   usr_rx3_pma_pll_lock_track_o   : out std_logic
);
end NX_HSSL_U_FULL;
--#}}}#

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_HSSL_U_FULL definition                                                           2019/06/20
-- =================================================================================================

-- NX_HSSL_U_FULL#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

architecture NX_RTL of NX_HSSL_U_FULL is

signal LINK_RX0 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX1 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX2 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_RX3 : std_logic_vector(CRX_LINK_SIZE-1 downto 0);
signal LINK_TX0 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX1 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX2 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);
signal LINK_TX3 : std_logic_vector(CTX_LINK_SIZE-1 downto 0);

-- component NX_CTX_U#{{{#
component NX_CTX_U
 generic (
     cfg_tx_pcs_protocol_size_i    : bit := '0';
     cfg_tx_pcs_8b_scr_sel_i       : bit := '0';
     cfg_tx_pcs_scr_init_i         : bit_vector(16 downto 0) := (others => '0');
     cfg_tx_pcs_scr_bypass_i       : bit := '0';
     cfg_tx_pcs_sync_supported_i   : bit := '0';
     cfg_tx_pcs_replace_bypass_i   : bit := '0';
     cfg_tx_pcs_enc_bypass_i       : bit := '0';
     cfg_tx_pcs_loopback_i         : bit := '0';
     cfg_tx_pcs_polarity_i         : bit := '0';
     cfg_tx_pcs_esistream_fsm_en_i : bit := '0';
     cfg_tx_pcs_bypass_pma_cdc_i   : bit := '0';
     cfg_tx_pcs_bypass_usr_cdc_i   : bit := '0';
     cfg_tx_pma_clk_pos_i          : bit := '0';
     cfg_tx_pma_loopback_i         : bit := '0';
     cfg_tx_gearbox_en_i           : bit := '0';
     cfg_tx_gearbox_mode_i         : bit := '0';

     location             : string := ""
 );
port (
    ENC_E_I1 : in  std_logic;
    ENC_E_I2 : in  std_logic;
    ENC_E_I3 : in  std_logic;
    ENC_E_I4 : in  std_logic;
    ENC_E_I5 : in  std_logic;
    ENC_E_I6 : in  std_logic;
    ENC_E_I7 : in  std_logic;
    ENC_E_I8 : in  std_logic;

    CH_K_I1  : in  std_logic;
    CH_K_I2  : in  std_logic;
    CH_K_I3  : in  std_logic;
    CH_K_I4  : in  std_logic;
    CH_K_I5  : in  std_logic;
    CH_K_I6  : in  std_logic;
    CH_K_I7  : in  std_logic;
    CH_K_I8  : in  std_logic;

    SCR_E_I1 : in  std_logic;
    SCR_E_I2 : in  std_logic;
    SCR_E_I3 : in  std_logic;
    SCR_E_I4 : in  std_logic;
    SCR_E_I5 : in  std_logic;
    SCR_E_I6 : in  std_logic;
    SCR_E_I7 : in  std_logic;
    SCR_E_I8 : in  std_logic;

    EOMF_I1  : in  std_logic;
    EOMF_I2  : in  std_logic;
    EOMF_I3  : in  std_logic;
    EOMF_I4  : in  std_logic;
    EOMF_I5  : in  std_logic;
    EOMF_I6  : in  std_logic;
    EOMF_I7  : in  std_logic;
    EOMF_I8  : in  std_logic;

    EOF_I1   : in  std_logic;
    EOF_I2   : in  std_logic;
    EOF_I3   : in  std_logic;
    EOF_I4   : in  std_logic;
    EOF_I5   : in  std_logic;
    EOF_I6   : in  std_logic;
    EOF_I7   : in  std_logic;
    EOF_I8   : in  std_logic;

    REP_E_I  : in  std_logic;
    RST_N_I  : in  std_logic;

    PWDN_N_I : in  std_logic;

    DATA_I1  : in  std_logic;
    DATA_I2  : in  std_logic;
    DATA_I3  : in  std_logic;
    DATA_I4  : in  std_logic;
    DATA_I5  : in  std_logic;
    DATA_I6  : in  std_logic;
    DATA_I7  : in  std_logic;
    DATA_I8  : in  std_logic;
    DATA_I9  : in  std_logic;
    DATA_I10 : in  std_logic;
    DATA_I11 : in  std_logic;
    DATA_I12 : in  std_logic;
    DATA_I13 : in  std_logic;
    DATA_I14 : in  std_logic;
    DATA_I15 : in  std_logic;
    DATA_I16 : in  std_logic;
    DATA_I17 : in  std_logic;
    DATA_I18 : in  std_logic;
    DATA_I19 : in  std_logic;
    DATA_I20 : in  std_logic;
    DATA_I21 : in  std_logic;
    DATA_I22 : in  std_logic;
    DATA_I23 : in  std_logic;
    DATA_I24 : in  std_logic;
    DATA_I25 : in  std_logic;
    DATA_I26 : in  std_logic;
    DATA_I27 : in  std_logic;
    DATA_I28 : in  std_logic;
    DATA_I29 : in  std_logic;
    DATA_I30 : in  std_logic;
    DATA_I31 : in  std_logic;
    DATA_I32 : in  std_logic;
    DATA_I33 : in  std_logic;
    DATA_I34 : in  std_logic;
    DATA_I35 : in  std_logic;
    DATA_I36 : in  std_logic;
    DATA_I37 : in  std_logic;
    DATA_I38 : in  std_logic;
    DATA_I39 : in  std_logic;
    DATA_I40 : in  std_logic;
    DATA_I41 : in  std_logic;
    DATA_I42 : in  std_logic;
    DATA_I43 : in  std_logic;
    DATA_I44 : in  std_logic;
    DATA_I45 : in  std_logic;
    DATA_I46 : in  std_logic;
    DATA_I47 : in  std_logic;
    DATA_I48 : in  std_logic;
    DATA_I49 : in  std_logic;
    DATA_I50 : in  std_logic;
    DATA_I51 : in  std_logic;
    DATA_I52 : in  std_logic;
    DATA_I53 : in  std_logic;
    DATA_I54 : in  std_logic;
    DATA_I55 : in  std_logic;
    DATA_I56 : in  std_logic;
    DATA_I57 : in  std_logic;
    DATA_I58 : in  std_logic;
    DATA_I59 : in  std_logic;
    DATA_I60 : in  std_logic;
    DATA_I61 : in  std_logic;
    DATA_I62 : in  std_logic;
    DATA_I63 : in  std_logic;
    DATA_I64 : in  std_logic;

    INV_K_O  : out std_logic;
    CLK_O    : out std_logic;

    BUSY_O   : out std_logic;
    CLK_E_I  : in  std_logic;


    LINK     : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0)
);
end component;
--#}}}#

-- component NX_CRX_U#{{{#
component NX_CRX_U
 generic (
     cfg_rx_pma_m_eye_ppm_i                     : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_coarse_ppm_i                    : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_fine_ppm_i                      : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_cmd_i               : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_peak_detect_on_i                : bit := '0';
     cfg_rx_pma_dco_reg_res_i                   : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_vref_sel_i                  : bit := '0';
     cfg_rx_pma_dco_divl_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_dco_divm_i                      : bit := '0';
     cfg_rx_pma_dco_divn_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_loopback_i                      : bit := '0';
     cfg_rx_pma_clk_pos_i                       : bit := '0';
     cfg_rx_pma_cdr_cp_i                        : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pma_ctrl_term_i                     : bit_vector(5 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divm_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_divn_en_n_i                 : bit := '0';
     cfg_rx_pma_pll_cpump_n_i                   : bit_vector(2 downto 0) := (others => '0');
     cfg_rx_pma_pll_divf_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divm_i                      : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pma_pll_divn_i                      : bit := '0';
     cfg_rx_pcs_debug_en_i                      : bit := '0';
     cfg_rx_pcs_bypass_pma_cdc_i                : bit := '0';
     cfg_rx_pcs_fsm_watchdog_en_i               : bit := '0';
     cfg_rx_pcs_fsm_sel_i                       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_polarity_i                      : bit := '0';
     cfg_rx_pcs_loopback_i                      : bit := '0';
     cfg_rx_pcs_dscr_bypass_i                   : bit := '0';
     cfg_rx_pcs_8b_dscr_sel_i                   : bit := '0';
     cfg_rx_pcs_replace_bypass_i                : bit := '0';
     cfg_rx_pcs_sync_supported_i                : bit := '0';
     cfg_rx_pcs_buffers_bypass_i                : bit := '0';
     cfg_rx_pcs_buffers_use_cdc_i               : bit := '0';
     cfg_rx_pcs_el_buff_skp_header_3_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_2_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_1_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_0_i          : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_header_size_i       : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_3_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_2_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_1_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_char_0_i            : bit_vector(8 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_skp_seq_size_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_only_one_skp_i          : bit := '0';
     cfg_rx_pcs_el_buff_diff_bef_comp_i         : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_el_buff_max_comp_i              : bit_vector(3 downto 0) := (others => '0');
     cfg_rx_pcs_dec_bypass_i                    : bit := '0';
     cfg_rx_pcs_align_bypass_i                  : bit := '0';
     cfg_rx_pcs_nb_comma_bef_realign_i          : bit_vector(1 downto 0) := (others => '0');
     cfg_rx_pcs_comma_mask_i                    : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_m_comma_en_i                    : bit := '0';
     cfg_rx_pcs_p_comma_val_i                   : bit_vector(9 downto 0) := (others => '0');
     cfg_rx_pcs_p_comma_en_i                    : bit := '0';
     cfg_rx_pcs_bypass_usr_cdc_i                : bit := '0';
     cfg_rx_pcs_protocol_size_i                 : bit := '0';
     cfg_rx_gearbox_mode_i                      : bit := '0';
     cfg_rx_gearbox_en_i                        : bit := '0';

     location                     : string := ""
 );
port (
    DSCR_E_I  : in  std_logic;
    DEC_E_I   : in  std_logic;
    ALIGN_E_I : in  std_logic;
    ALIGN_S_I : in  std_logic;
    REP_E_I   : in  std_logic;
    BUF_R_I   : in  std_logic;

    OVS_BS_I1 : in  std_logic;
    OVS_BS_I2 : in  std_logic;

    RST_N_I   : in  std_logic;

    PMA_RSTN_I: in  std_logic;
    MEYE_RST_I: in  std_logic;
    PWDN_N_I  : in  std_logic;

    DBG_S_I1  : in  std_logic;
    DBG_S_I2  : in  std_logic;
    DBG_S_I3  : in  std_logic;

    DATA_O1   : out std_logic;
    DATA_O2   : out std_logic;
    DATA_O3   : out std_logic;
    DATA_O4   : out std_logic;
    DATA_O5   : out std_logic;
    DATA_O6   : out std_logic;
    DATA_O7   : out std_logic;
    DATA_O8   : out std_logic;
    DATA_O9   : out std_logic;
    DATA_O10  : out std_logic;
    DATA_O11  : out std_logic;
    DATA_O12  : out std_logic;
    DATA_O13  : out std_logic;
    DATA_O14  : out std_logic;
    DATA_O15  : out std_logic;
    DATA_O16  : out std_logic;
    DATA_O17  : out std_logic;
    DATA_O18  : out std_logic;
    DATA_O19  : out std_logic;
    DATA_O20  : out std_logic;
    DATA_O21  : out std_logic;
    DATA_O22  : out std_logic;
    DATA_O23  : out std_logic;
    DATA_O24  : out std_logic;
    DATA_O25  : out std_logic;
    DATA_O26  : out std_logic;
    DATA_O27  : out std_logic;
    DATA_O28  : out std_logic;
    DATA_O29  : out std_logic;
    DATA_O30  : out std_logic;
    DATA_O31  : out std_logic;
    DATA_O32  : out std_logic;
    DATA_O33  : out std_logic;
    DATA_O34  : out std_logic;
    DATA_O35  : out std_logic;
    DATA_O36  : out std_logic;
    DATA_O37  : out std_logic;
    DATA_O38  : out std_logic;
    DATA_O39  : out std_logic;
    DATA_O40  : out std_logic;
    DATA_O41  : out std_logic;
    DATA_O42  : out std_logic;
    DATA_O43  : out std_logic;
    DATA_O44  : out std_logic;
    DATA_O45  : out std_logic;
    DATA_O46  : out std_logic;
    DATA_O47  : out std_logic;
    DATA_O48  : out std_logic;
    DATA_O49  : out std_logic;
    DATA_O50  : out std_logic;
    DATA_O51  : out std_logic;
    DATA_O52  : out std_logic;
    DATA_O53  : out std_logic;
    DATA_O54  : out std_logic;
    DATA_O55  : out std_logic;
    DATA_O56  : out std_logic;
    DATA_O57  : out std_logic;
    DATA_O58  : out std_logic;
    DATA_O59  : out std_logic;
    DATA_O60  : out std_logic;
    DATA_O61  : out std_logic;
    DATA_O62  : out std_logic;
    DATA_O63  : out std_logic;
    DATA_O64  : out std_logic;

    CH_COM_O1 : out std_logic;
    CH_COM_O2 : out std_logic;
    CH_COM_O3 : out std_logic;
    CH_COM_O4 : out std_logic;
    CH_COM_O5 : out std_logic;
    CH_COM_O6 : out std_logic;
    CH_COM_O7 : out std_logic;
    CH_COM_O8 : out std_logic;

    CH_K_O1   : out std_logic;
    CH_K_O2   : out std_logic;
    CH_K_O3   : out std_logic;
    CH_K_O4   : out std_logic;
    CH_K_O5   : out std_logic;
    CH_K_O6   : out std_logic;
    CH_K_O7   : out std_logic;
    CH_K_O8   : out std_logic;

    NIT_O1    : out std_logic;
    NIT_O2    : out std_logic;
    NIT_O3    : out std_logic;
    NIT_O4    : out std_logic;
    NIT_O5    : out std_logic;
    NIT_O6    : out std_logic;
    NIT_O7    : out std_logic;
    NIT_O8    : out std_logic;

    D_ERR_O1  : out std_logic;
    D_ERR_O2  : out std_logic;
    D_ERR_O3  : out std_logic;
    D_ERR_O4  : out std_logic;
    D_ERR_O5  : out std_logic;
    D_ERR_O6  : out std_logic;
    D_ERR_O7  : out std_logic;
    D_ERR_O8  : out std_logic;

    CH_A_O1   : out std_logic;
    CH_A_O2   : out std_logic;
    CH_A_O3   : out std_logic;
    CH_A_O4   : out std_logic;
    CH_A_O5   : out std_logic;
    CH_A_O6   : out std_logic;
    CH_A_O7   : out std_logic;
    CH_A_O8   : out std_logic;

    CH_F_O1   : out std_logic;
    CH_F_O2   : out std_logic;
    CH_F_O3   : out std_logic;
    CH_F_O4   : out std_logic;
    CH_F_O5   : out std_logic;
    CH_F_O6   : out std_logic;
    CH_F_O7   : out std_logic;
    CH_F_O8   : out std_logic;

    ALIGN_O    : out std_logic;
    VREALIGN_O : out std_logic;
    BUSY_O     : out std_logic;

    TST_O1    : out std_logic;
    TST_O2    : out std_logic;
    TST_O3    : out std_logic;
    TST_O4    : out std_logic;
    TST_O5    : out std_logic;
    TST_O6    : out std_logic;
    TST_O7    : out std_logic;
    TST_O8    : out std_logic;

    LOS_O     : out std_logic;

    LL_FLOCK_O  : out std_logic;
    LL_SLOCK_O  : out std_logic;
    PLL_LOCK_O  : out std_logic;
    PLL_LOCKT_O : out std_logic;

    LINK      : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0)
);
end component;
--#}}}#

-- component NX_PMA_U#{{{#
component NX_PMA_U
generic (
   cfg_pll_pma_int_data_len_i            : bit := '0';
   cfg_pll_pma_cpump_i                   : bit_vector( 3 downto 0) := (others => '0');
   cfg_pll_pma_divl_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_divm_i                    : bit := '0';
   cfg_pll_pma_divn_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_lvds_en_i                 : bit := '0';
   cfg_pll_pma_lvds_mux_i                : bit := '0';
   cfg_pll_pma_mux_ckref_i               : bit := '0';
   cfg_pll_pma_gbx_en_i                  : bit := '0';
   cfg_pll_pma_ckref_ext_i               : bit := '0';
   cfg_main_clk_to_fabric_div_mode_i     : bit := '0';
   cfg_main_clk_to_fabric_div_en_i       : bit := '0';
   cfg_main_clk_to_fabric_sel_i          : bit := '0';
   cfg_main_rclk_to_fabric_sel_i         : bit_vector( 1 downto 0) := (others => '0');
   cfg_main_use_only_usr_clock_i         : bit := '0';
   tx_usrclk_use_pcs_clk_2               : bit := '0';
   rx_usrclk_use_pcs_clk_2               : bit := '0';
   cfg_pcs_word_len_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pcs_ovs_en_i                      : bit := '0';
   cfg_pcs_ovs_mode_i                    : bit := '0';
   cfg_pcs_pll_lock_ppm_i                : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_m_eye_i            : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_up_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_dn_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_coarse_ena_i : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_fine_ena_i   : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_step_i       : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_mode_i        : bit_vector( 1 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_locked_i      : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_unlocked_i    : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_1        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_2        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx1_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx2_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx3_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx0_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx1_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx2_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx3_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx0_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_test_mode_i                       : bit_vector( 1 downto 0) := (others => '0');

   location                    : string := ""
);
port (
    CLK_TX_I    : in  std_logic;
    CLK_RX_I    : in  std_logic;
    CLK_REF_I   : in  std_logic;

    DC_E_I       : in  std_logic;
    DC_LCSN_I1   : in  std_logic;
    DC_LCSN_I2   : in  std_logic;
    DC_LCSN_I3   : in  std_logic;
    DC_LCSN_I4   : in  std_logic;

    DC_CCSN_I    : in  std_logic;
    DC_WE_N_I    : in  std_logic;

    DC_ADD_I1    : in  std_logic;
    DC_ADD_I2    : in  std_logic;
    DC_ADD_I3    : in  std_logic;
    DC_ADD_I4    : in  std_logic;
    DC_WDATAS_I  : in  std_logic;
    DC_WDATA_I1  : in  std_logic;
    DC_WDATA_I2  : in  std_logic;
    DC_WDATA_I3  : in  std_logic;
    DC_WDATA_I4  : in  std_logic;
    DC_WDATA_I5  : in  std_logic;
    DC_WDATA_I6  : in  std_logic;
    DC_WDATA_I7  : in  std_logic;
    DC_WDATA_I8  : in  std_logic;
    DC_WDATA_I9  : in  std_logic;
    DC_WDATA_I10 : in  std_logic;
    DC_WDATA_I11 : in  std_logic;
    DC_WDATA_I12 : in  std_logic;

    PLL_RN_I     : in  std_logic;
    PWDN_N_I     : in  std_logic;
    RST_N_I      : in  std_logic;

    DBG_S_I1     : in  std_logic;
    DBG_S_I2     : in  std_logic;
    DBG_A_I      : in  std_logic;

    SE_I         : in  std_logic;

    SCAN_I1      : in  std_logic;
    SCAN_I2      : in  std_logic;
    SCAN_I3      : in  std_logic;
    SCAN_I4      : in  std_logic;
    SCAN_I5      : in  std_logic;
    SCAN_I6      : in  std_logic;
    SCAN_I7      : in  std_logic;
    SCAN_I8      : in  std_logic;

    CLK_O       : out std_logic;
    CLK_RX_O    : out std_logic;
    LOCK_O      : out std_logic;
    LOCKA_O     : out std_logic;
    FB_LOCK_O   : out std_logic;
    CAL_OUT_O   : out std_logic;
    DBG_R_O     : out std_logic;

    LL_O1       : out std_logic;
    LL_O2       : out std_logic;
    LL_O3       : out std_logic;
    LL_O4       : out std_logic;
    LL_O5       : out std_logic;
    LL_O6       : out std_logic;
    LL_O7       : out std_logic;
    LL_O8       : out std_logic;
    LL_O9       : out std_logic;
    LL_O10      : out std_logic;
    LL_O11      : out std_logic;
    LL_O12      : out std_logic;
    LL_O13      : out std_logic;
    LL_O14      : out std_logic;
    LL_O15      : out std_logic;
    LL_O16      : out std_logic;
    LL_O17      : out std_logic;
    LL_O18      : out std_logic;
    LL_O19      : out std_logic;
    LL_O20      : out std_logic;


    SCAN_O1     : out std_logic;
    SCAN_O2     : out std_logic;
    SCAN_O3     : out std_logic;
    SCAN_O4     : out std_logic;
    SCAN_O5     : out std_logic;
    SCAN_O6     : out std_logic;
    SCAN_O7     : out std_logic;
    SCAN_O8     : out std_logic;


    LINK_TX0    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX1    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX2    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX3    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_RX0    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX1    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX2    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX3    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0)
);
end component;
--#}}}#

begin

-- ctrl: NX_PMA_U#{{{#
ctrl: NX_PMA_U generic map (
    cfg_pll_pma_int_data_len_i              => cfg_pll_pma_int_data_len_i
  , cfg_pll_pma_cpump_i                     => cfg_pll_pma_cpump_i
  , cfg_pll_pma_divl_i                      => cfg_pll_pma_divl_i
  , cfg_pll_pma_divm_i                      => cfg_pll_pma_divm_i
  , cfg_pll_pma_divn_i                      => cfg_pll_pma_divn_i
  , cfg_pll_pma_lvds_en_i                   => cfg_pll_pma_lvds_en_i
  , cfg_pll_pma_lvds_mux_i                  => cfg_pll_pma_lvds_mux_i
  , cfg_pll_pma_mux_ckref_i                 => cfg_pll_pma_mux_ckref_i
  , cfg_pll_pma_gbx_en_i                    => cfg_pll_pma_gbx_en_i
  , cfg_pll_pma_ckref_ext_i                 => cfg_pll_pma_ckref_ext_i
  , cfg_main_clk_to_fabric_div_mode_i       => cfg_main_clk_to_fabric_div_mode_i
  , cfg_main_clk_to_fabric_div_en_i         => cfg_main_clk_to_fabric_div_en_i
  , cfg_main_clk_to_fabric_sel_i            => cfg_main_clk_to_fabric_sel_i
  , cfg_main_rclk_to_fabric_sel_i           => cfg_main_rclk_to_fabric_sel_i
  , cfg_main_use_only_usr_clock_i           => cfg_main_use_only_usr_clock_i
  , tx_usrclk_use_pcs_clk_2                 => tx_usrclk_use_pcs_clk_2
  , rx_usrclk_use_pcs_clk_2                 => rx_usrclk_use_pcs_clk_2
  , cfg_pcs_word_len_i                      => cfg_pcs_word_len_i
  , cfg_pcs_ovs_en_i                        => cfg_pcs_ovs_en_i
  , cfg_pcs_ovs_mode_i                      => cfg_pcs_ovs_mode_i
  , cfg_pcs_pll_lock_ppm_i                  => cfg_pcs_pll_lock_ppm_i
  , cfg_dyn_all_rx_pma_m_eye_i              => cfg_dyn_all_rx_pma_m_eye_i
  , cfg_dyn_all_rx_pma_m_eye_up_i           => cfg_dyn_all_rx_pma_m_eye_up_i
  , cfg_dyn_all_rx_pma_m_eye_dn_i           => cfg_dyn_all_rx_pma_m_eye_dn_i
  , cfg_dyn_all_rx_pma_m_eye_coarse_ena_i   => cfg_dyn_all_rx_pma_m_eye_coarse_ena_i
  , cfg_dyn_all_rx_pma_m_eye_fine_ena_i     => cfg_dyn_all_rx_pma_m_eye_fine_ena_i
  , cfg_dyn_all_rx_pma_m_eye_step_i         => cfg_dyn_all_rx_pma_m_eye_step_i
  , cfg_dyn_all_rx_pma_trim_mode_i          => cfg_dyn_all_rx_pma_trim_mode_i
  , cfg_dyn_all_rx_pma_trim_locked_i        => cfg_dyn_all_rx_pma_trim_locked_i
  , cfg_dyn_all_rx_pma_trim_unlocked_i      => cfg_dyn_all_rx_pma_trim_unlocked_i
  , cfg_dyn_all_rx_pma_threshold_1          => cfg_dyn_all_rx_pma_threshold_1
  , cfg_dyn_all_rx_pma_threshold_2          => cfg_dyn_all_rx_pma_threshold_2
  , cfg_dyn_tx0_pma_pre_sign_i              => cfg_dyn_tx0_pma_pre_sign_i
  , cfg_dyn_tx1_pma_pre_sign_i              => cfg_dyn_tx1_pma_pre_sign_i
  , cfg_dyn_tx2_pma_pre_sign_i              => cfg_dyn_tx2_pma_pre_sign_i
  , cfg_dyn_tx3_pma_pre_sign_i              => cfg_dyn_tx3_pma_pre_sign_i
  , cfg_dyn_tx0_pma_pre_en_i                => cfg_dyn_tx0_pma_pre_en_i
  , cfg_dyn_tx1_pma_pre_en_i                => cfg_dyn_tx1_pma_pre_en_i
  , cfg_dyn_tx2_pma_pre_en_i                => cfg_dyn_tx2_pma_pre_en_i
  , cfg_dyn_tx3_pma_pre_en_i                => cfg_dyn_tx3_pma_pre_en_i
  , cfg_dyn_tx0_pma_pre_sel_i               => cfg_dyn_tx0_pma_pre_sel_i
  , cfg_dyn_tx1_pma_pre_sel_i               => cfg_dyn_tx1_pma_pre_sel_i
  , cfg_dyn_tx2_pma_pre_sel_i               => cfg_dyn_tx2_pma_pre_sel_i
  , cfg_dyn_tx3_pma_pre_sel_i               => cfg_dyn_tx3_pma_pre_sel_i
  , cfg_dyn_tx0_pma_main_sign_i             => cfg_dyn_tx0_pma_main_sign_i
  , cfg_dyn_tx1_pma_main_sign_i             => cfg_dyn_tx1_pma_main_sign_i
  , cfg_dyn_tx2_pma_main_sign_i             => cfg_dyn_tx2_pma_main_sign_i
  , cfg_dyn_tx3_pma_main_sign_i             => cfg_dyn_tx3_pma_main_sign_i
  , cfg_dyn_tx0_pma_main_en_i               => cfg_dyn_tx0_pma_main_en_i
  , cfg_dyn_tx1_pma_main_en_i               => cfg_dyn_tx1_pma_main_en_i
  , cfg_dyn_tx2_pma_main_en_i               => cfg_dyn_tx2_pma_main_en_i
  , cfg_dyn_tx3_pma_main_en_i               => cfg_dyn_tx3_pma_main_en_i
  , cfg_dyn_tx0_pma_margin_sel_i            => cfg_dyn_tx0_pma_margin_sel_i
  , cfg_dyn_tx1_pma_margin_sel_i            => cfg_dyn_tx1_pma_margin_sel_i
  , cfg_dyn_tx2_pma_margin_sel_i            => cfg_dyn_tx2_pma_margin_sel_i
  , cfg_dyn_tx3_pma_margin_sel_i            => cfg_dyn_tx3_pma_margin_sel_i
  , cfg_dyn_tx0_pma_margin_input_i          => cfg_dyn_tx0_pma_margin_input_i
  , cfg_dyn_tx1_pma_margin_input_i          => cfg_dyn_tx1_pma_margin_input_i
  , cfg_dyn_tx2_pma_margin_input_i          => cfg_dyn_tx2_pma_margin_input_i
  , cfg_dyn_tx3_pma_margin_input_i          => cfg_dyn_tx3_pma_margin_input_i
  , cfg_dyn_tx0_pma_post_sign_i             => cfg_dyn_tx0_pma_post_sign_i
  , cfg_dyn_tx1_pma_post_sign_i             => cfg_dyn_tx1_pma_post_sign_i
  , cfg_dyn_tx2_pma_post_sign_i             => cfg_dyn_tx2_pma_post_sign_i
  , cfg_dyn_tx3_pma_post_sign_i             => cfg_dyn_tx3_pma_post_sign_i
  , cfg_dyn_tx0_pma_post_en_i               => cfg_dyn_tx0_pma_post_en_i
  , cfg_dyn_tx1_pma_post_en_i               => cfg_dyn_tx1_pma_post_en_i
  , cfg_dyn_tx2_pma_post_en_i               => cfg_dyn_tx2_pma_post_en_i
  , cfg_dyn_tx3_pma_post_en_i               => cfg_dyn_tx3_pma_post_en_i
  , cfg_dyn_tx0_pma_post_sel_i              => cfg_dyn_tx0_pma_post_sel_i
  , cfg_dyn_tx1_pma_post_sel_i              => cfg_dyn_tx1_pma_post_sel_i
  , cfg_dyn_tx2_pma_post_sel_i              => cfg_dyn_tx2_pma_post_sel_i
  , cfg_dyn_tx3_pma_post_sel_i              => cfg_dyn_tx3_pma_post_sel_i
  , cfg_dyn_rx0_pma_ctle_cap_p_i            => cfg_dyn_rx0_pma_ctle_cap_p_i
  , cfg_dyn_rx1_pma_ctle_cap_p_i            => cfg_dyn_rx1_pma_ctle_cap_p_i
  , cfg_dyn_rx2_pma_ctle_cap_p_i            => cfg_dyn_rx2_pma_ctle_cap_p_i
  , cfg_dyn_rx3_pma_ctle_cap_p_i            => cfg_dyn_rx3_pma_ctle_cap_p_i
  , cfg_dyn_rx0_pma_ctle_res_p_i            => cfg_dyn_rx0_pma_ctle_res_p_i
  , cfg_dyn_rx1_pma_ctle_res_p_i            => cfg_dyn_rx1_pma_ctle_res_p_i
  , cfg_dyn_rx2_pma_ctle_res_p_i            => cfg_dyn_rx2_pma_ctle_res_p_i
  , cfg_dyn_rx3_pma_ctle_res_p_i            => cfg_dyn_rx3_pma_ctle_res_p_i
  , cfg_dyn_rx0_pma_dfe_idac_tap1_n_i       => cfg_dyn_rx0_pma_dfe_idac_tap1_n_i
  , cfg_dyn_rx1_pma_dfe_idac_tap1_n_i       => cfg_dyn_rx1_pma_dfe_idac_tap1_n_i
  , cfg_dyn_rx2_pma_dfe_idac_tap1_n_i       => cfg_dyn_rx2_pma_dfe_idac_tap1_n_i
  , cfg_dyn_rx3_pma_dfe_idac_tap1_n_i       => cfg_dyn_rx3_pma_dfe_idac_tap1_n_i
  , cfg_dyn_rx0_pma_dfe_idac_tap2_n_i       => cfg_dyn_rx0_pma_dfe_idac_tap2_n_i
  , cfg_dyn_rx1_pma_dfe_idac_tap2_n_i       => cfg_dyn_rx1_pma_dfe_idac_tap2_n_i
  , cfg_dyn_rx2_pma_dfe_idac_tap2_n_i       => cfg_dyn_rx2_pma_dfe_idac_tap2_n_i
  , cfg_dyn_rx3_pma_dfe_idac_tap2_n_i       => cfg_dyn_rx3_pma_dfe_idac_tap2_n_i
  , cfg_dyn_rx0_pma_dfe_idac_tap3_n_i       => cfg_dyn_rx0_pma_dfe_idac_tap3_n_i
  , cfg_dyn_rx1_pma_dfe_idac_tap3_n_i       => cfg_dyn_rx1_pma_dfe_idac_tap3_n_i
  , cfg_dyn_rx2_pma_dfe_idac_tap3_n_i       => cfg_dyn_rx2_pma_dfe_idac_tap3_n_i
  , cfg_dyn_rx3_pma_dfe_idac_tap3_n_i       => cfg_dyn_rx3_pma_dfe_idac_tap3_n_i
  , cfg_dyn_rx0_pma_dfe_idac_tap4_n_i       => cfg_dyn_rx0_pma_dfe_idac_tap4_n_i
  , cfg_dyn_rx1_pma_dfe_idac_tap4_n_i       => cfg_dyn_rx1_pma_dfe_idac_tap4_n_i
  , cfg_dyn_rx2_pma_dfe_idac_tap4_n_i       => cfg_dyn_rx2_pma_dfe_idac_tap4_n_i
  , cfg_dyn_rx3_pma_dfe_idac_tap4_n_i       => cfg_dyn_rx3_pma_dfe_idac_tap4_n_i
  , cfg_dyn_rx0_pma_termination_cmd_i       => cfg_dyn_rx0_pma_termination_cmd_i
  , cfg_dyn_rx1_pma_termination_cmd_i       => cfg_dyn_rx1_pma_termination_cmd_i
  , cfg_dyn_rx2_pma_termination_cmd_i       => cfg_dyn_rx2_pma_termination_cmd_i
  , cfg_dyn_rx3_pma_termination_cmd_i       => cfg_dyn_rx3_pma_termination_cmd_i
  , cfg_test_mode_i                         => cfg_test_mode_i

  , location                                => location & ":COMMON1.PMA1"
 )
port map (
    CLK_TX_I       => hssl_clk_user_tx_i
  , CLK_RX_I       => hssl_clk_user_rx_i
  , CLK_REF_I      => hssl_clk_ref_i
  , CLK_O          => hssl_clock_o
  , CLK_RX_O       => hssl_rclock_o
  , DC_E_I         => usr_dyn_cfg_en_i
  , DC_LCSN_I1     => usr_dyn_cfg_lane_cs_n_i(0)
  , DC_LCSN_I2     => usr_dyn_cfg_lane_cs_n_i(1)
  , DC_LCSN_I3     => usr_dyn_cfg_lane_cs_n_i(2)
  , DC_LCSN_I4     => usr_dyn_cfg_lane_cs_n_i(3)
  , DC_CCSN_I      => usr_dyn_cfg_calibration_cs_n_i
  , DC_WE_N_I      => usr_dyn_cfg_we_n_i
  , DC_ADD_I1      => usr_dyn_cfg_addr_i(0)
  , DC_ADD_I2      => usr_dyn_cfg_addr_i(1)
  , DC_ADD_I3      => usr_dyn_cfg_addr_i(2)
  , DC_ADD_I4      => usr_dyn_cfg_addr_i(3)
  , DC_WDATAS_I    => usr_dyn_cfg_wdata_sel_i
  , DC_WDATA_I1    => usr_dyn_cfg_wdata_i(0)
  , DC_WDATA_I2    => usr_dyn_cfg_wdata_i(1)
  , DC_WDATA_I3    => usr_dyn_cfg_wdata_i(2)
  , DC_WDATA_I4    => usr_dyn_cfg_wdata_i(3)
  , DC_WDATA_I5    => usr_dyn_cfg_wdata_i(4)
  , DC_WDATA_I6    => usr_dyn_cfg_wdata_i(5)
  , DC_WDATA_I7    => usr_dyn_cfg_wdata_i(6)
  , DC_WDATA_I8    => usr_dyn_cfg_wdata_i(7)
  , DC_WDATA_I9    => usr_dyn_cfg_wdata_i(8)
  , DC_WDATA_I10   => usr_dyn_cfg_wdata_i(9)
  , DC_WDATA_I11   => usr_dyn_cfg_wdata_i(10)
  , DC_WDATA_I12   => usr_dyn_cfg_wdata_i(11)
  , PLL_RN_I       => usr_pll_pma_rst_n_i
  , PWDN_N_I       => usr_pll_pma_pwr_down_n_i
  , RST_N_I        => usr_main_rst_n_i
  , LOCK_O         => usr_pll_lock_o
  , LOCKA_O        => usr_pll_pma_lock_analog_o
  , FB_LOCK_O      => usr_pll_ckfb_lock_o
  , CAL_OUT_O      => usr_calibrate_pma_out_o
  , DBG_S_I1       => usr_main_async_debug_lane_sel_i(0)
  , DBG_S_I2       => usr_main_async_debug_lane_sel_i(1)
  , DBG_A_I        => usr_main_async_debug_ack_i
  , DBG_R_O        => usr_main_async_debug_req_o
  , LL_O1          => usr_main_rx_pma_ll_out_o(0)
  , LL_O2          => usr_main_rx_pma_ll_out_o(1)
  , LL_O3          => usr_main_rx_pma_ll_out_o(2)
  , LL_O4          => usr_main_rx_pma_ll_out_o(3)
  , LL_O5          => usr_main_rx_pma_ll_out_o(4)
  , LL_O6          => usr_main_rx_pma_ll_out_o(5)
  , LL_O7          => usr_main_rx_pma_ll_out_o(6)
  , LL_O8          => usr_main_rx_pma_ll_out_o(7)
  , LL_O9          => usr_main_rx_pma_ll_out_o(8)
  , LL_O10         => usr_main_rx_pma_ll_out_o(9)
  , LL_O11         => usr_main_rx_pma_ll_out_o(10)
  , LL_O12         => usr_main_rx_pma_ll_out_o(11)
  , LL_O13         => usr_main_rx_pma_ll_out_o(12)
  , LL_O14         => usr_main_rx_pma_ll_out_o(13)
  , LL_O15         => usr_main_rx_pma_ll_out_o(14)
  , LL_O16         => usr_main_rx_pma_ll_out_o(15)
  , LL_O17         => usr_main_rx_pma_ll_out_o(16)
  , LL_O18         => usr_main_rx_pma_ll_out_o(17)
  , LL_O19         => usr_main_rx_pma_ll_out_o(18)
  , LL_O20         => usr_main_rx_pma_ll_out_o(19)
  , SE_I           => scan_en_i
  , SCAN_I1        => scan_in_i(0)
  , SCAN_I2        => scan_in_i(1)
  , SCAN_I3        => scan_in_i(2)
  , SCAN_I4        => scan_in_i(3)
  , SCAN_I5        => scan_in_i(4)
  , SCAN_I6        => scan_in_i(5)
  , SCAN_I7        => scan_in_i(6)
  , SCAN_I8        => scan_in_i(7)
  , SCAN_O1        => scan_out_o(0)
  , SCAN_O2        => scan_out_o(1)
  , SCAN_O3        => scan_out_o(2)
  , SCAN_O4        => scan_out_o(3)
  , SCAN_O5        => scan_out_o(4)
  , SCAN_O6        => scan_out_o(5)
  , SCAN_O7        => scan_out_o(6)
  , SCAN_O8        => scan_out_o(7)

  , LINK_TX0       => LINK_TX0
  , LINK_TX1       => LINK_TX1
  , LINK_TX2       => LINK_TX2
  , LINK_TX3       => LINK_TX3
  , LINK_RX0       => LINK_RX0
  , LINK_RX1       => LINK_RX1
  , LINK_RX2       => LINK_RX2
  , LINK_RX3       => LINK_RX3
);
--#}}}#

-- txlane0: NX_CTX_U#{{{#
txlane0: NX_CTX_U generic map (
   cfg_tx_pcs_protocol_size_i    => cfg_tx0_pcs_protocol_size_i
 , cfg_tx_pcs_8b_scr_sel_i       => cfg_tx0_pcs_8b_scr_sel_i
 , cfg_tx_pcs_scr_init_i         => cfg_tx0_pcs_scr_init_i
 , cfg_tx_pcs_scr_bypass_i       => cfg_tx0_pcs_scr_bypass_i
 , cfg_tx_pcs_sync_supported_i   => cfg_tx0_pcs_sync_supported_i
 , cfg_tx_pcs_replace_bypass_i   => cfg_tx0_pcs_replace_bypass_i
 , cfg_tx_pcs_enc_bypass_i       => cfg_tx0_pcs_enc_bypass_i
 , cfg_tx_pcs_loopback_i         => cfg_tx0_pcs_loopback_i
 , cfg_tx_pcs_polarity_i         => cfg_tx0_pcs_polarity_i
 , cfg_tx_pcs_esistream_fsm_en_i => cfg_tx0_pcs_esistream_fsm_en_i
 , cfg_tx_pcs_bypass_pma_cdc_i   => cfg_tx0_pcs_bypass_pma_cdc_i
 , cfg_tx_pcs_bypass_usr_cdc_i   => cfg_tx0_pcs_bypass_usr_cdc_i
 , cfg_tx_pma_clk_pos_i          => cfg_tx0_pma_clk_pos_i
 , cfg_tx_pma_loopback_i         => cfg_tx0_pma_loopback_i
 , cfg_tx_gearbox_en_i           => cfg_tx0_gearbox_en_i
 , cfg_tx_gearbox_mode_i         => cfg_tx0_gearbox_mode_i
 , location                      => location & ":CHANNEL1.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx0_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx0_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx0_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx0_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx0_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx0_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx0_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx0_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx0_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx0_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx0_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx0_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx0_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx0_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx0_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx0_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx0_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx0_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx0_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx0_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx0_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx0_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx0_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx0_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx0_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx0_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx0_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx0_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx0_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx0_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx0_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx0_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx0_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx0_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx0_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx0_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx0_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx0_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx0_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx0_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx0_ctrl_replace_en_i
  , RST_N_I  => usr_tx0_rst_n_i

  , DATA_I1  => usr_tx0_data_i(0)
  , DATA_I2  => usr_tx0_data_i(1)
  , DATA_I3  => usr_tx0_data_i(2)
  , DATA_I4  => usr_tx0_data_i(3)
  , DATA_I5  => usr_tx0_data_i(4)
  , DATA_I6  => usr_tx0_data_i(5)
  , DATA_I7  => usr_tx0_data_i(6)
  , DATA_I8  => usr_tx0_data_i(7)
  , DATA_I9  => usr_tx0_data_i(8)
  , DATA_I10 => usr_tx0_data_i(9)
  , DATA_I11 => usr_tx0_data_i(10)
  , DATA_I12 => usr_tx0_data_i(11)
  , DATA_I13 => usr_tx0_data_i(12)
  , DATA_I14 => usr_tx0_data_i(13)
  , DATA_I15 => usr_tx0_data_i(14)
  , DATA_I16 => usr_tx0_data_i(15)
  , DATA_I17 => usr_tx0_data_i(16)
  , DATA_I18 => usr_tx0_data_i(17)
  , DATA_I19 => usr_tx0_data_i(18)
  , DATA_I20 => usr_tx0_data_i(19)
  , DATA_I21 => usr_tx0_data_i(20)
  , DATA_I22 => usr_tx0_data_i(21)
  , DATA_I23 => usr_tx0_data_i(22)
  , DATA_I24 => usr_tx0_data_i(23)
  , DATA_I25 => usr_tx0_data_i(24)
  , DATA_I26 => usr_tx0_data_i(25)
  , DATA_I27 => usr_tx0_data_i(26)
  , DATA_I28 => usr_tx0_data_i(27)
  , DATA_I29 => usr_tx0_data_i(28)
  , DATA_I30 => usr_tx0_data_i(29)
  , DATA_I31 => usr_tx0_data_i(30)
  , DATA_I32 => usr_tx0_data_i(31)
  , DATA_I33 => usr_tx0_data_i(32)
  , DATA_I34 => usr_tx0_data_i(33)
  , DATA_I35 => usr_tx0_data_i(34)
  , DATA_I36 => usr_tx0_data_i(35)
  , DATA_I37 => usr_tx0_data_i(36)
  , DATA_I38 => usr_tx0_data_i(37)
  , DATA_I39 => usr_tx0_data_i(38)
  , DATA_I40 => usr_tx0_data_i(39)
  , DATA_I41 => usr_tx0_data_i(40)
  , DATA_I42 => usr_tx0_data_i(41)
  , DATA_I43 => usr_tx0_data_i(42)
  , DATA_I44 => usr_tx0_data_i(43)
  , DATA_I45 => usr_tx0_data_i(44)
  , DATA_I46 => usr_tx0_data_i(45)
  , DATA_I47 => usr_tx0_data_i(46)
  , DATA_I48 => usr_tx0_data_i(47)
  , DATA_I49 => usr_tx0_data_i(48)
  , DATA_I50 => usr_tx0_data_i(49)
  , DATA_I51 => usr_tx0_data_i(50)
  , DATA_I52 => usr_tx0_data_i(51)
  , DATA_I53 => usr_tx0_data_i(52)
  , DATA_I54 => usr_tx0_data_i(53)
  , DATA_I55 => usr_tx0_data_i(54)
  , DATA_I56 => usr_tx0_data_i(55)
  , DATA_I57 => usr_tx0_data_i(56)
  , DATA_I58 => usr_tx0_data_i(57)
  , DATA_I59 => usr_tx0_data_i(58)
  , DATA_I60 => usr_tx0_data_i(59)
  , DATA_I61 => usr_tx0_data_i(60)
  , DATA_I62 => usr_tx0_data_i(61)
  , DATA_I63 => usr_tx0_data_i(62)
  , DATA_I64 => usr_tx0_data_i(63)

  , BUSY_O   => usr_tx0_busy_o
  , INV_K_O  => usr_tx0_ctrl_invalid_k_o

  , PWDN_N_I => usr_tx0_ctrl_driver_pwrdwn_n_i
  , CLK_E_I  => usr_tx0_pma_clk_en_i
  , CLK_O    => usr_tx0_pma_tx_clk_o

  , LINK     => LINK_TX0
);
--#}}}#

-- rxlane0: NX_CRX_U#{{{#
rxlane0: NX_CRX_U generic map (
    cfg_rx_pma_m_eye_ppm_i               => cfg_rx0_pma_m_eye_ppm_i
  , cfg_rx_pma_coarse_ppm_i              => cfg_rx0_pma_coarse_ppm_i
  , cfg_rx_pma_fine_ppm_i                => cfg_rx0_pma_fine_ppm_i
  , cfg_rx_pma_peak_detect_cmd_i         => cfg_rx0_pma_peak_detect_cmd_i
  , cfg_rx_pma_peak_detect_on_i          => cfg_rx0_pma_peak_detect_on_i
  , cfg_rx_pma_dco_reg_res_i             => cfg_rx0_pma_dco_reg_res_i
  , cfg_rx_pma_dco_vref_sel_i            => cfg_rx0_pma_dco_vref_sel_i
  , cfg_rx_pma_dco_divl_i                => cfg_rx0_pma_dco_divl_i
  , cfg_rx_pma_dco_divm_i                => cfg_rx0_pma_dco_divm_i
  , cfg_rx_pma_dco_divn_i                => cfg_rx0_pma_dco_divn_i
  , cfg_rx_pma_loopback_i                => cfg_rx0_pma_loopback_i
  , cfg_rx_pma_clk_pos_i                 => cfg_rx0_pma_clk_pos_i
  , cfg_rx_pma_cdr_cp_i                  => cfg_rx0_pma_cdr_cp_i
  , cfg_rx_pma_ctrl_term_i               => cfg_rx0_pma_ctrl_term_i
  , cfg_rx_pma_pll_divf_en_n_i           => cfg_rx0_pma_pll_divf_en_n_i
  , cfg_rx_pma_pll_divm_en_n_i           => cfg_rx0_pma_pll_divm_en_n_i
  , cfg_rx_pma_pll_divn_en_n_i           => cfg_rx0_pma_pll_divn_en_n_i
  , cfg_rx_pma_pll_cpump_n_i             => cfg_rx0_pma_pll_cpump_n_i
  , cfg_rx_pma_pll_divf_i                => cfg_rx0_pma_pll_divf_i
  , cfg_rx_pma_pll_divm_i                => cfg_rx0_pma_pll_divm_i
  , cfg_rx_pma_pll_divn_i                => cfg_rx0_pma_pll_divn_i
  , cfg_rx_pcs_debug_en_i                => cfg_rx0_pcs_debug_en_i
  , cfg_rx_pcs_bypass_pma_cdc_i          => cfg_rx0_pcs_bypass_pma_cdc_i
  , cfg_rx_pcs_fsm_watchdog_en_i         => cfg_rx0_pcs_fsm_watchdog_en_i
  , cfg_rx_pcs_fsm_sel_i                 => cfg_rx0_pcs_fsm_sel_i
  , cfg_rx_pcs_polarity_i                => cfg_rx0_pcs_polarity_i
  , cfg_rx_pcs_loopback_i                => cfg_rx0_pcs_loopback_i
  , cfg_rx_pcs_dscr_bypass_i             => cfg_rx0_pcs_dscr_bypass_i
  , cfg_rx_pcs_8b_dscr_sel_i             => cfg_rx0_pcs_8b_dscr_sel_i
  , cfg_rx_pcs_replace_bypass_i          => cfg_rx0_pcs_replace_bypass_i
  , cfg_rx_pcs_sync_supported_i          => cfg_rx0_pcs_sync_supported_i
  , cfg_rx_pcs_buffers_bypass_i          => cfg_rx0_pcs_buffers_bypass_i
  , cfg_rx_pcs_buffers_use_cdc_i         => cfg_rx0_pcs_buffers_use_cdc_i
  , cfg_rx_pcs_el_buff_skp_header_3_i    => cfg_rx0_pcs_el_buff_skp_header_3_i
  , cfg_rx_pcs_el_buff_skp_header_2_i    => cfg_rx0_pcs_el_buff_skp_header_2_i
  , cfg_rx_pcs_el_buff_skp_header_1_i    => cfg_rx0_pcs_el_buff_skp_header_1_i
  , cfg_rx_pcs_el_buff_skp_header_0_i    => cfg_rx0_pcs_el_buff_skp_header_0_i
  , cfg_rx_pcs_el_buff_skp_header_size_i => cfg_rx0_pcs_el_buff_skp_header_size_i
  , cfg_rx_pcs_el_buff_skp_char_3_i      => cfg_rx0_pcs_el_buff_skp_char_3_i
  , cfg_rx_pcs_el_buff_skp_char_2_i      => cfg_rx0_pcs_el_buff_skp_char_2_i
  , cfg_rx_pcs_el_buff_skp_char_1_i      => cfg_rx0_pcs_el_buff_skp_char_1_i
  , cfg_rx_pcs_el_buff_skp_char_0_i      => cfg_rx0_pcs_el_buff_skp_char_0_i
  , cfg_rx_pcs_el_buff_skp_seq_size_i    => cfg_rx0_pcs_el_buff_skp_seq_size_i
  , cfg_rx_pcs_el_buff_only_one_skp_i    => cfg_rx0_pcs_el_buff_only_one_skp_i
  , cfg_rx_pcs_el_buff_diff_bef_comp_i   => cfg_rx0_pcs_el_buff_diff_bef_comp_i
  , cfg_rx_pcs_el_buff_max_comp_i        => cfg_rx0_pcs_el_buff_max_comp_i
  , cfg_rx_pcs_dec_bypass_i              => cfg_rx0_pcs_dec_bypass_i
  , cfg_rx_pcs_align_bypass_i            => cfg_rx0_pcs_align_bypass_i
  , cfg_rx_pcs_nb_comma_bef_realign_i    => cfg_rx0_pcs_nb_comma_bef_realign_i
  , cfg_rx_pcs_comma_mask_i              => cfg_rx0_pcs_comma_mask_i
  , cfg_rx_pcs_m_comma_val_i             => cfg_rx0_pcs_m_comma_val_i
  , cfg_rx_pcs_m_comma_en_i              => cfg_rx0_pcs_m_comma_en_i
  , cfg_rx_pcs_p_comma_val_i             => cfg_rx0_pcs_p_comma_val_i
  , cfg_rx_pcs_p_comma_en_i              => cfg_rx0_pcs_p_comma_en_i
  , cfg_rx_pcs_bypass_usr_cdc_i          => cfg_rx0_pcs_bypass_usr_cdc_i
  , cfg_rx_pcs_protocol_size_i           => cfg_rx0_pcs_protocol_size_i
  , cfg_rx_gearbox_mode_i                => cfg_rx0_gearbox_mode_i
  , cfg_rx_gearbox_en_i                  => cfg_rx0_gearbox_en_i
  , location                             => location & ":CHANNEL1.CRX1"
 )
port map (
    DSCR_E_I    => usr_rx0_ctrl_dscr_en_i
  , DEC_E_I     => usr_rx0_ctrl_dec_en_i
  , ALIGN_E_I   => usr_rx0_ctrl_align_en_i
  , ALIGN_S_I   => usr_rx0_ctrl_align_sync_i
  , REP_E_I     => usr_rx0_ctrl_replace_en_i
  , BUF_R_I     => usr_rx0_ctrl_el_buff_rst_i

  , OVS_BS_I1   => usr_rx0_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2   => usr_rx0_ctrl_ovs_bit_sel_i(1)

  , RST_N_I     => usr_rx0_rst_n_i

  , PMA_RSTN_I  => usr_rx0_pma_rst_n_i
  , MEYE_RST_I  => usr_rx0_pma_m_eye_rst_i
  , PWDN_N_I    => usr_rx0_pma_pwr_down_n_i
  , DBG_S_I1    => usr_rx0_ctrl_debug_sel_i(0)
  , DBG_S_I2    => usr_rx0_ctrl_debug_sel_i(1)
  , DBG_S_I3    => usr_rx0_ctrl_debug_sel_i(2)

  , DATA_O1     => usr_rx0_data_o(0)
  , DATA_O2     => usr_rx0_data_o(1)
  , DATA_O3     => usr_rx0_data_o(2)
  , DATA_O4     => usr_rx0_data_o(3)
  , DATA_O5     => usr_rx0_data_o(4)
  , DATA_O6     => usr_rx0_data_o(5)
  , DATA_O7     => usr_rx0_data_o(6)
  , DATA_O8     => usr_rx0_data_o(7)
  , DATA_O9     => usr_rx0_data_o(8)
  , DATA_O10    => usr_rx0_data_o(9)
  , DATA_O11    => usr_rx0_data_o(10)
  , DATA_O12    => usr_rx0_data_o(11)
  , DATA_O13    => usr_rx0_data_o(12)
  , DATA_O14    => usr_rx0_data_o(13)
  , DATA_O15    => usr_rx0_data_o(14)
  , DATA_O16    => usr_rx0_data_o(15)
  , DATA_O17    => usr_rx0_data_o(16)
  , DATA_O18    => usr_rx0_data_o(17)
  , DATA_O19    => usr_rx0_data_o(18)
  , DATA_O20    => usr_rx0_data_o(19)
  , DATA_O21    => usr_rx0_data_o(20)
  , DATA_O22    => usr_rx0_data_o(21)
  , DATA_O23    => usr_rx0_data_o(22)
  , DATA_O24    => usr_rx0_data_o(23)
  , DATA_O25    => usr_rx0_data_o(24)
  , DATA_O26    => usr_rx0_data_o(25)
  , DATA_O27    => usr_rx0_data_o(26)
  , DATA_O28    => usr_rx0_data_o(27)
  , DATA_O29    => usr_rx0_data_o(28)
  , DATA_O30    => usr_rx0_data_o(29)
  , DATA_O31    => usr_rx0_data_o(30)
  , DATA_O32    => usr_rx0_data_o(31)
  , DATA_O33    => usr_rx0_data_o(32)
  , DATA_O34    => usr_rx0_data_o(33)
  , DATA_O35    => usr_rx0_data_o(34)
  , DATA_O36    => usr_rx0_data_o(35)
  , DATA_O37    => usr_rx0_data_o(36)
  , DATA_O38    => usr_rx0_data_o(37)
  , DATA_O39    => usr_rx0_data_o(38)
  , DATA_O40    => usr_rx0_data_o(39)
  , DATA_O41    => usr_rx0_data_o(40)
  , DATA_O42    => usr_rx0_data_o(41)
  , DATA_O43    => usr_rx0_data_o(42)
  , DATA_O44    => usr_rx0_data_o(43)
  , DATA_O45    => usr_rx0_data_o(44)
  , DATA_O46    => usr_rx0_data_o(45)
  , DATA_O47    => usr_rx0_data_o(46)
  , DATA_O48    => usr_rx0_data_o(47)
  , DATA_O49    => usr_rx0_data_o(48)
  , DATA_O50    => usr_rx0_data_o(49)
  , DATA_O51    => usr_rx0_data_o(50)
  , DATA_O52    => usr_rx0_data_o(51)
  , DATA_O53    => usr_rx0_data_o(52)
  , DATA_O54    => usr_rx0_data_o(53)
  , DATA_O55    => usr_rx0_data_o(54)
  , DATA_O56    => usr_rx0_data_o(55)
  , DATA_O57    => usr_rx0_data_o(56)
  , DATA_O58    => usr_rx0_data_o(57)
  , DATA_O59    => usr_rx0_data_o(58)
  , DATA_O60    => usr_rx0_data_o(59)
  , DATA_O61    => usr_rx0_data_o(60)
  , DATA_O62    => usr_rx0_data_o(61)
  , DATA_O63    => usr_rx0_data_o(62)
  , DATA_O64    => usr_rx0_data_o(63)

  , CH_COM_O1   => usr_rx0_ctrl_char_is_comma_o(0)
  , CH_COM_O2   => usr_rx0_ctrl_char_is_comma_o(1)
  , CH_COM_O3   => usr_rx0_ctrl_char_is_comma_o(2)
  , CH_COM_O4   => usr_rx0_ctrl_char_is_comma_o(3)
  , CH_COM_O5   => usr_rx0_ctrl_char_is_comma_o(4)
  , CH_COM_O6   => usr_rx0_ctrl_char_is_comma_o(5)
  , CH_COM_O7   => usr_rx0_ctrl_char_is_comma_o(6)
  , CH_COM_O8   => usr_rx0_ctrl_char_is_comma_o(7)

  , CH_K_O1     => usr_rx0_ctrl_char_is_k_o(0)
  , CH_K_O2     => usr_rx0_ctrl_char_is_k_o(1)
  , CH_K_O3     => usr_rx0_ctrl_char_is_k_o(2)
  , CH_K_O4     => usr_rx0_ctrl_char_is_k_o(3)
  , CH_K_O5     => usr_rx0_ctrl_char_is_k_o(4)
  , CH_K_O6     => usr_rx0_ctrl_char_is_k_o(5)
  , CH_K_O7     => usr_rx0_ctrl_char_is_k_o(6)
  , CH_K_O8     => usr_rx0_ctrl_char_is_k_o(7)

  , NIT_O1      => usr_rx0_ctrl_not_in_table_o(0)
  , NIT_O2      => usr_rx0_ctrl_not_in_table_o(1)
  , NIT_O3      => usr_rx0_ctrl_not_in_table_o(2)
  , NIT_O4      => usr_rx0_ctrl_not_in_table_o(3)
  , NIT_O5      => usr_rx0_ctrl_not_in_table_o(4)
  , NIT_O6      => usr_rx0_ctrl_not_in_table_o(5)
  , NIT_O7      => usr_rx0_ctrl_not_in_table_o(6)
  , NIT_O8      => usr_rx0_ctrl_not_in_table_o(7)

  , D_ERR_O1    => usr_rx0_ctrl_disp_err_o(0)
  , D_ERR_O2    => usr_rx0_ctrl_disp_err_o(1)
  , D_ERR_O3    => usr_rx0_ctrl_disp_err_o(2)
  , D_ERR_O4    => usr_rx0_ctrl_disp_err_o(3)
  , D_ERR_O5    => usr_rx0_ctrl_disp_err_o(4)
  , D_ERR_O6    => usr_rx0_ctrl_disp_err_o(5)
  , D_ERR_O7    => usr_rx0_ctrl_disp_err_o(6)
  , D_ERR_O8    => usr_rx0_ctrl_disp_err_o(7)

  , CH_A_O1     => usr_rx0_ctrl_char_is_a_o(0)
  , CH_A_O2     => usr_rx0_ctrl_char_is_a_o(1)
  , CH_A_O3     => usr_rx0_ctrl_char_is_a_o(2)
  , CH_A_O4     => usr_rx0_ctrl_char_is_a_o(3)
  , CH_A_O5     => usr_rx0_ctrl_char_is_a_o(4)
  , CH_A_O6     => usr_rx0_ctrl_char_is_a_o(5)
  , CH_A_O7     => usr_rx0_ctrl_char_is_a_o(6)
  , CH_A_O8     => usr_rx0_ctrl_char_is_a_o(7)

  , CH_F_O1     => usr_rx0_ctrl_char_is_f_o(0)
  , CH_F_O2     => usr_rx0_ctrl_char_is_f_o(1)
  , CH_F_O3     => usr_rx0_ctrl_char_is_f_o(2)
  , CH_F_O4     => usr_rx0_ctrl_char_is_f_o(3)
  , CH_F_O5     => usr_rx0_ctrl_char_is_f_o(4)
  , CH_F_O6     => usr_rx0_ctrl_char_is_f_o(5)
  , CH_F_O7     => usr_rx0_ctrl_char_is_f_o(6)
  , CH_F_O8     => usr_rx0_ctrl_char_is_f_o(7)

  , ALIGN_O     => usr_rx0_ctrl_char_is_aligned_o
  , VREALIGN_O  => usr_rx0_ctrl_valid_realign_o
  , BUSY_O      => usr_rx0_busy_o

  , TST_O1      => usr_rx0_test_o(0)
  , TST_O2      => usr_rx0_test_o(1)
  , TST_O3      => usr_rx0_test_o(2)
  , TST_O4      => usr_rx0_test_o(3)
  , TST_O5      => usr_rx0_test_o(4)
  , TST_O6      => usr_rx0_test_o(5)
  , TST_O7      => usr_rx0_test_o(6)
  , TST_O8      => usr_rx0_test_o(7)

  , LOS_O       => usr_rx0_pma_loss_of_signal_o
  , LL_FLOCK_O  => usr_rx0_pma_ll_fast_locked_o
  , LL_SLOCK_O  => usr_rx0_pma_ll_slow_locked_o
  , PLL_LOCK_O  => usr_rx0_pma_pll_lock_o
  , PLL_LOCKT_O => usr_rx0_pma_pll_lock_track_o

  , LINK       => LINK_RX0
);
--#}}}#

-- txlane1: NX_CTX_U#{{{#
txlane1: NX_CTX_U generic map (

   cfg_tx_pcs_protocol_size_i    => cfg_tx1_pcs_protocol_size_i
 , cfg_tx_pcs_8b_scr_sel_i       => cfg_tx1_pcs_8b_scr_sel_i
 , cfg_tx_pcs_scr_init_i         => cfg_tx1_pcs_scr_init_i
 , cfg_tx_pcs_scr_bypass_i       => cfg_tx1_pcs_scr_bypass_i
 , cfg_tx_pcs_sync_supported_i   => cfg_tx1_pcs_sync_supported_i
 , cfg_tx_pcs_replace_bypass_i   => cfg_tx1_pcs_replace_bypass_i
 , cfg_tx_pcs_enc_bypass_i       => cfg_tx1_pcs_enc_bypass_i
 , cfg_tx_pcs_loopback_i         => cfg_tx1_pcs_loopback_i
 , cfg_tx_pcs_polarity_i         => cfg_tx1_pcs_polarity_i
 , cfg_tx_pcs_esistream_fsm_en_i => cfg_tx1_pcs_esistream_fsm_en_i
 , cfg_tx_pcs_bypass_pma_cdc_i   => cfg_tx1_pcs_bypass_pma_cdc_i
 , cfg_tx_pcs_bypass_usr_cdc_i   => cfg_tx1_pcs_bypass_usr_cdc_i
 , cfg_tx_pma_clk_pos_i          => cfg_tx1_pma_clk_pos_i
 , cfg_tx_pma_loopback_i         => cfg_tx1_pma_loopback_i
 , cfg_tx_gearbox_en_i           => cfg_tx1_gearbox_en_i
 , cfg_tx_gearbox_mode_i         => cfg_tx1_gearbox_mode_i
 , location                      => location & ":CHANNEL2.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx1_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx1_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx1_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx1_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx1_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx1_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx1_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx1_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx1_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx1_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx1_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx1_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx1_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx1_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx1_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx1_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx1_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx1_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx1_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx1_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx1_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx1_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx1_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx1_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx1_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx1_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx1_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx1_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx1_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx1_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx1_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx1_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx1_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx1_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx1_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx1_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx1_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx1_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx1_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx1_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx1_ctrl_replace_en_i
  , RST_N_I  => usr_tx1_rst_n_i

  , DATA_I1  => usr_tx1_data_i(0)
  , DATA_I2  => usr_tx1_data_i(1)
  , DATA_I3  => usr_tx1_data_i(2)
  , DATA_I4  => usr_tx1_data_i(3)
  , DATA_I5  => usr_tx1_data_i(4)
  , DATA_I6  => usr_tx1_data_i(5)
  , DATA_I7  => usr_tx1_data_i(6)
  , DATA_I8  => usr_tx1_data_i(7)
  , DATA_I9  => usr_tx1_data_i(8)
  , DATA_I10 => usr_tx1_data_i(9)
  , DATA_I11 => usr_tx1_data_i(10)
  , DATA_I12 => usr_tx1_data_i(11)
  , DATA_I13 => usr_tx1_data_i(12)
  , DATA_I14 => usr_tx1_data_i(13)
  , DATA_I15 => usr_tx1_data_i(14)
  , DATA_I16 => usr_tx1_data_i(15)
  , DATA_I17 => usr_tx1_data_i(16)
  , DATA_I18 => usr_tx1_data_i(17)
  , DATA_I19 => usr_tx1_data_i(18)
  , DATA_I20 => usr_tx1_data_i(19)
  , DATA_I21 => usr_tx1_data_i(20)
  , DATA_I22 => usr_tx1_data_i(21)
  , DATA_I23 => usr_tx1_data_i(22)
  , DATA_I24 => usr_tx1_data_i(23)
  , DATA_I25 => usr_tx1_data_i(24)
  , DATA_I26 => usr_tx1_data_i(25)
  , DATA_I27 => usr_tx1_data_i(26)
  , DATA_I28 => usr_tx1_data_i(27)
  , DATA_I29 => usr_tx1_data_i(28)
  , DATA_I30 => usr_tx1_data_i(29)
  , DATA_I31 => usr_tx1_data_i(30)
  , DATA_I32 => usr_tx1_data_i(31)
  , DATA_I33 => usr_tx1_data_i(32)
  , DATA_I34 => usr_tx1_data_i(33)
  , DATA_I35 => usr_tx1_data_i(34)
  , DATA_I36 => usr_tx1_data_i(35)
  , DATA_I37 => usr_tx1_data_i(36)
  , DATA_I38 => usr_tx1_data_i(37)
  , DATA_I39 => usr_tx1_data_i(38)
  , DATA_I40 => usr_tx1_data_i(39)
  , DATA_I41 => usr_tx1_data_i(40)
  , DATA_I42 => usr_tx1_data_i(41)
  , DATA_I43 => usr_tx1_data_i(42)
  , DATA_I44 => usr_tx1_data_i(43)
  , DATA_I45 => usr_tx1_data_i(44)
  , DATA_I46 => usr_tx1_data_i(45)
  , DATA_I47 => usr_tx1_data_i(46)
  , DATA_I48 => usr_tx1_data_i(47)
  , DATA_I49 => usr_tx1_data_i(48)
  , DATA_I50 => usr_tx1_data_i(49)
  , DATA_I51 => usr_tx1_data_i(50)
  , DATA_I52 => usr_tx1_data_i(51)
  , DATA_I53 => usr_tx1_data_i(52)
  , DATA_I54 => usr_tx1_data_i(53)
  , DATA_I55 => usr_tx1_data_i(54)
  , DATA_I56 => usr_tx1_data_i(55)
  , DATA_I57 => usr_tx1_data_i(56)
  , DATA_I58 => usr_tx1_data_i(57)
  , DATA_I59 => usr_tx1_data_i(58)
  , DATA_I60 => usr_tx1_data_i(59)
  , DATA_I61 => usr_tx1_data_i(60)
  , DATA_I62 => usr_tx1_data_i(61)
  , DATA_I63 => usr_tx1_data_i(62)
  , DATA_I64 => usr_tx1_data_i(63)

  , BUSY_O   => usr_tx1_busy_o
  , INV_K_O  => usr_tx1_ctrl_invalid_k_o

  , PWDN_N_I => usr_tx1_ctrl_driver_pwrdwn_n_i
  , CLK_E_I  => usr_tx1_pma_clk_en_i
  , CLK_O    => usr_tx1_pma_tx_clk_o

  , LINK     => LINK_TX1
);
--#}}}#

-- rxlane1: NX_CRX_U#{{{#
rxlane1: NX_CRX_U generic map (
    cfg_rx_pma_m_eye_ppm_i               => cfg_rx1_pma_m_eye_ppm_i
  , cfg_rx_pma_coarse_ppm_i              => cfg_rx1_pma_coarse_ppm_i
  , cfg_rx_pma_fine_ppm_i                => cfg_rx1_pma_fine_ppm_i
  , cfg_rx_pma_peak_detect_cmd_i         => cfg_rx1_pma_peak_detect_cmd_i
  , cfg_rx_pma_peak_detect_on_i          => cfg_rx1_pma_peak_detect_on_i
  , cfg_rx_pma_dco_reg_res_i             => cfg_rx1_pma_dco_reg_res_i
  , cfg_rx_pma_dco_vref_sel_i            => cfg_rx1_pma_dco_vref_sel_i
  , cfg_rx_pma_dco_divl_i                => cfg_rx1_pma_dco_divl_i
  , cfg_rx_pma_dco_divm_i                => cfg_rx1_pma_dco_divm_i
  , cfg_rx_pma_dco_divn_i                => cfg_rx1_pma_dco_divn_i
  , cfg_rx_pma_loopback_i                => cfg_rx1_pma_loopback_i
  , cfg_rx_pma_clk_pos_i                 => cfg_rx1_pma_clk_pos_i
  , cfg_rx_pma_cdr_cp_i                  => cfg_rx1_pma_cdr_cp_i
  , cfg_rx_pma_ctrl_term_i               => cfg_rx1_pma_ctrl_term_i
  , cfg_rx_pma_pll_divf_en_n_i           => cfg_rx1_pma_pll_divf_en_n_i
  , cfg_rx_pma_pll_divm_en_n_i           => cfg_rx1_pma_pll_divm_en_n_i
  , cfg_rx_pma_pll_divn_en_n_i           => cfg_rx1_pma_pll_divn_en_n_i
  , cfg_rx_pma_pll_cpump_n_i             => cfg_rx1_pma_pll_cpump_n_i
  , cfg_rx_pma_pll_divf_i                => cfg_rx1_pma_pll_divf_i
  , cfg_rx_pma_pll_divm_i                => cfg_rx1_pma_pll_divm_i
  , cfg_rx_pma_pll_divn_i                => cfg_rx1_pma_pll_divn_i
  , cfg_rx_pcs_debug_en_i                => cfg_rx1_pcs_debug_en_i
  , cfg_rx_pcs_bypass_pma_cdc_i          => cfg_rx1_pcs_bypass_pma_cdc_i
  , cfg_rx_pcs_fsm_watchdog_en_i         => cfg_rx1_pcs_fsm_watchdog_en_i
  , cfg_rx_pcs_fsm_sel_i                 => cfg_rx1_pcs_fsm_sel_i
  , cfg_rx_pcs_polarity_i                => cfg_rx1_pcs_polarity_i
  , cfg_rx_pcs_loopback_i                => cfg_rx1_pcs_loopback_i
  , cfg_rx_pcs_dscr_bypass_i             => cfg_rx1_pcs_dscr_bypass_i
  , cfg_rx_pcs_8b_dscr_sel_i             => cfg_rx1_pcs_8b_dscr_sel_i
  , cfg_rx_pcs_replace_bypass_i          => cfg_rx1_pcs_replace_bypass_i
  , cfg_rx_pcs_sync_supported_i          => cfg_rx1_pcs_sync_supported_i
  , cfg_rx_pcs_buffers_bypass_i          => cfg_rx1_pcs_buffers_bypass_i
  , cfg_rx_pcs_buffers_use_cdc_i         => cfg_rx1_pcs_buffers_use_cdc_i
  , cfg_rx_pcs_el_buff_skp_header_3_i    => cfg_rx1_pcs_el_buff_skp_header_3_i
  , cfg_rx_pcs_el_buff_skp_header_2_i    => cfg_rx1_pcs_el_buff_skp_header_2_i
  , cfg_rx_pcs_el_buff_skp_header_1_i    => cfg_rx1_pcs_el_buff_skp_header_1_i
  , cfg_rx_pcs_el_buff_skp_header_0_i    => cfg_rx1_pcs_el_buff_skp_header_0_i
  , cfg_rx_pcs_el_buff_skp_header_size_i => cfg_rx1_pcs_el_buff_skp_header_size_i
  , cfg_rx_pcs_el_buff_skp_char_3_i      => cfg_rx1_pcs_el_buff_skp_char_3_i
  , cfg_rx_pcs_el_buff_skp_char_2_i      => cfg_rx1_pcs_el_buff_skp_char_2_i
  , cfg_rx_pcs_el_buff_skp_char_1_i      => cfg_rx1_pcs_el_buff_skp_char_1_i
  , cfg_rx_pcs_el_buff_skp_char_0_i      => cfg_rx1_pcs_el_buff_skp_char_0_i
  , cfg_rx_pcs_el_buff_skp_seq_size_i    => cfg_rx1_pcs_el_buff_skp_seq_size_i
  , cfg_rx_pcs_el_buff_only_one_skp_i    => cfg_rx1_pcs_el_buff_only_one_skp_i
  , cfg_rx_pcs_el_buff_diff_bef_comp_i   => cfg_rx1_pcs_el_buff_diff_bef_comp_i
  , cfg_rx_pcs_el_buff_max_comp_i        => cfg_rx1_pcs_el_buff_max_comp_i
  , cfg_rx_pcs_dec_bypass_i              => cfg_rx1_pcs_dec_bypass_i
  , cfg_rx_pcs_align_bypass_i            => cfg_rx1_pcs_align_bypass_i
  , cfg_rx_pcs_nb_comma_bef_realign_i    => cfg_rx1_pcs_nb_comma_bef_realign_i
  , cfg_rx_pcs_comma_mask_i              => cfg_rx1_pcs_comma_mask_i
  , cfg_rx_pcs_m_comma_val_i             => cfg_rx1_pcs_m_comma_val_i
  , cfg_rx_pcs_m_comma_en_i              => cfg_rx1_pcs_m_comma_en_i
  , cfg_rx_pcs_p_comma_val_i             => cfg_rx1_pcs_p_comma_val_i
  , cfg_rx_pcs_p_comma_en_i              => cfg_rx1_pcs_p_comma_en_i
  , cfg_rx_pcs_bypass_usr_cdc_i          => cfg_rx1_pcs_bypass_usr_cdc_i
  , cfg_rx_pcs_protocol_size_i           => cfg_rx1_pcs_protocol_size_i
  , cfg_rx_gearbox_mode_i                => cfg_rx1_gearbox_mode_i
  , cfg_rx_gearbox_en_i                  => cfg_rx1_gearbox_en_i
  , location                             => location & ":CHANNEL2.CRX1"
 )
port map (
    DSCR_E_I    => usr_rx1_ctrl_dscr_en_i
  , DEC_E_I     => usr_rx1_ctrl_dec_en_i
  , ALIGN_E_I   => usr_rx1_ctrl_align_en_i
  , ALIGN_S_I   => usr_rx1_ctrl_align_sync_i
  , REP_E_I     => usr_rx1_ctrl_replace_en_i
  , BUF_R_I     => usr_rx1_ctrl_el_buff_rst_i

  , OVS_BS_I1   => usr_rx1_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2   => usr_rx1_ctrl_ovs_bit_sel_i(1)

  , RST_N_I     => usr_rx1_rst_n_i

  , PMA_RSTN_I  => usr_rx1_pma_rst_n_i
  , MEYE_RST_I  => usr_rx1_pma_m_eye_rst_i
  , PWDN_N_I    => usr_rx1_pma_pwr_down_n_i
  , DBG_S_I1    => usr_rx1_ctrl_debug_sel_i(0)
  , DBG_S_I2    => usr_rx1_ctrl_debug_sel_i(1)
  , DBG_S_I3    => usr_rx1_ctrl_debug_sel_i(2)

  , DATA_O1     => usr_rx1_data_o(0)
  , DATA_O2     => usr_rx1_data_o(1)
  , DATA_O3     => usr_rx1_data_o(2)
  , DATA_O4     => usr_rx1_data_o(3)
  , DATA_O5     => usr_rx1_data_o(4)
  , DATA_O6     => usr_rx1_data_o(5)
  , DATA_O7     => usr_rx1_data_o(6)
  , DATA_O8     => usr_rx1_data_o(7)
  , DATA_O9     => usr_rx1_data_o(8)
  , DATA_O10    => usr_rx1_data_o(9)
  , DATA_O11    => usr_rx1_data_o(10)
  , DATA_O12    => usr_rx1_data_o(11)
  , DATA_O13    => usr_rx1_data_o(12)
  , DATA_O14    => usr_rx1_data_o(13)
  , DATA_O15    => usr_rx1_data_o(14)
  , DATA_O16    => usr_rx1_data_o(15)
  , DATA_O17    => usr_rx1_data_o(16)
  , DATA_O18    => usr_rx1_data_o(17)
  , DATA_O19    => usr_rx1_data_o(18)
  , DATA_O20    => usr_rx1_data_o(19)
  , DATA_O21    => usr_rx1_data_o(20)
  , DATA_O22    => usr_rx1_data_o(21)
  , DATA_O23    => usr_rx1_data_o(22)
  , DATA_O24    => usr_rx1_data_o(23)
  , DATA_O25    => usr_rx1_data_o(24)
  , DATA_O26    => usr_rx1_data_o(25)
  , DATA_O27    => usr_rx1_data_o(26)
  , DATA_O28    => usr_rx1_data_o(27)
  , DATA_O29    => usr_rx1_data_o(28)
  , DATA_O30    => usr_rx1_data_o(29)
  , DATA_O31    => usr_rx1_data_o(30)
  , DATA_O32    => usr_rx1_data_o(31)
  , DATA_O33    => usr_rx1_data_o(32)
  , DATA_O34    => usr_rx1_data_o(33)
  , DATA_O35    => usr_rx1_data_o(34)
  , DATA_O36    => usr_rx1_data_o(35)
  , DATA_O37    => usr_rx1_data_o(36)
  , DATA_O38    => usr_rx1_data_o(37)
  , DATA_O39    => usr_rx1_data_o(38)
  , DATA_O40    => usr_rx1_data_o(39)
  , DATA_O41    => usr_rx1_data_o(40)
  , DATA_O42    => usr_rx1_data_o(41)
  , DATA_O43    => usr_rx1_data_o(42)
  , DATA_O44    => usr_rx1_data_o(43)
  , DATA_O45    => usr_rx1_data_o(44)
  , DATA_O46    => usr_rx1_data_o(45)
  , DATA_O47    => usr_rx1_data_o(46)
  , DATA_O48    => usr_rx1_data_o(47)
  , DATA_O49    => usr_rx1_data_o(48)
  , DATA_O50    => usr_rx1_data_o(49)
  , DATA_O51    => usr_rx1_data_o(50)
  , DATA_O52    => usr_rx1_data_o(51)
  , DATA_O53    => usr_rx1_data_o(52)
  , DATA_O54    => usr_rx1_data_o(53)
  , DATA_O55    => usr_rx1_data_o(54)
  , DATA_O56    => usr_rx1_data_o(55)
  , DATA_O57    => usr_rx1_data_o(56)
  , DATA_O58    => usr_rx1_data_o(57)
  , DATA_O59    => usr_rx1_data_o(58)
  , DATA_O60    => usr_rx1_data_o(59)
  , DATA_O61    => usr_rx1_data_o(60)
  , DATA_O62    => usr_rx1_data_o(61)
  , DATA_O63    => usr_rx1_data_o(62)
  , DATA_O64    => usr_rx1_data_o(63)

  , CH_COM_O1   => usr_rx1_ctrl_char_is_comma_o(0)
  , CH_COM_O2   => usr_rx1_ctrl_char_is_comma_o(1)
  , CH_COM_O3   => usr_rx1_ctrl_char_is_comma_o(2)
  , CH_COM_O4   => usr_rx1_ctrl_char_is_comma_o(3)
  , CH_COM_O5   => usr_rx1_ctrl_char_is_comma_o(4)
  , CH_COM_O6   => usr_rx1_ctrl_char_is_comma_o(5)
  , CH_COM_O7   => usr_rx1_ctrl_char_is_comma_o(6)
  , CH_COM_O8   => usr_rx1_ctrl_char_is_comma_o(7)

  , CH_K_O1     => usr_rx1_ctrl_char_is_k_o(0)
  , CH_K_O2     => usr_rx1_ctrl_char_is_k_o(1)
  , CH_K_O3     => usr_rx1_ctrl_char_is_k_o(2)
  , CH_K_O4     => usr_rx1_ctrl_char_is_k_o(3)
  , CH_K_O5     => usr_rx1_ctrl_char_is_k_o(4)
  , CH_K_O6     => usr_rx1_ctrl_char_is_k_o(5)
  , CH_K_O7     => usr_rx1_ctrl_char_is_k_o(6)
  , CH_K_O8     => usr_rx1_ctrl_char_is_k_o(7)

  , NIT_O1      => usr_rx1_ctrl_not_in_table_o(0)
  , NIT_O2      => usr_rx1_ctrl_not_in_table_o(1)
  , NIT_O3      => usr_rx1_ctrl_not_in_table_o(2)
  , NIT_O4      => usr_rx1_ctrl_not_in_table_o(3)
  , NIT_O5      => usr_rx1_ctrl_not_in_table_o(4)
  , NIT_O6      => usr_rx1_ctrl_not_in_table_o(5)
  , NIT_O7      => usr_rx1_ctrl_not_in_table_o(6)
  , NIT_O8      => usr_rx1_ctrl_not_in_table_o(7)

  , D_ERR_O1    => usr_rx1_ctrl_disp_err_o(0)
  , D_ERR_O2    => usr_rx1_ctrl_disp_err_o(1)
  , D_ERR_O3    => usr_rx1_ctrl_disp_err_o(2)
  , D_ERR_O4    => usr_rx1_ctrl_disp_err_o(3)
  , D_ERR_O5    => usr_rx1_ctrl_disp_err_o(4)
  , D_ERR_O6    => usr_rx1_ctrl_disp_err_o(5)
  , D_ERR_O7    => usr_rx1_ctrl_disp_err_o(6)
  , D_ERR_O8    => usr_rx1_ctrl_disp_err_o(7)

  , CH_A_O1     => usr_rx1_ctrl_char_is_a_o(0)
  , CH_A_O2     => usr_rx1_ctrl_char_is_a_o(1)
  , CH_A_O3     => usr_rx1_ctrl_char_is_a_o(2)
  , CH_A_O4     => usr_rx1_ctrl_char_is_a_o(3)
  , CH_A_O5     => usr_rx1_ctrl_char_is_a_o(4)
  , CH_A_O6     => usr_rx1_ctrl_char_is_a_o(5)
  , CH_A_O7     => usr_rx1_ctrl_char_is_a_o(6)
  , CH_A_O8     => usr_rx1_ctrl_char_is_a_o(7)

  , CH_F_O1     => usr_rx1_ctrl_char_is_f_o(0)
  , CH_F_O2     => usr_rx1_ctrl_char_is_f_o(1)
  , CH_F_O3     => usr_rx1_ctrl_char_is_f_o(2)
  , CH_F_O4     => usr_rx1_ctrl_char_is_f_o(3)
  , CH_F_O5     => usr_rx1_ctrl_char_is_f_o(4)
  , CH_F_O6     => usr_rx1_ctrl_char_is_f_o(5)
  , CH_F_O7     => usr_rx1_ctrl_char_is_f_o(6)
  , CH_F_O8     => usr_rx1_ctrl_char_is_f_o(7)

  , ALIGN_O     => usr_rx1_ctrl_char_is_aligned_o
  , VREALIGN_O  => usr_rx1_ctrl_valid_realign_o
  , BUSY_O      => usr_rx1_busy_o

  , TST_O1      => usr_rx1_test_o(0)
  , TST_O2      => usr_rx1_test_o(1)
  , TST_O3      => usr_rx1_test_o(2)
  , TST_O4      => usr_rx1_test_o(3)
  , TST_O5      => usr_rx1_test_o(4)
  , TST_O6      => usr_rx1_test_o(5)
  , TST_O7      => usr_rx1_test_o(6)
  , TST_O8      => usr_rx1_test_o(7)

  , LOS_O       => usr_rx1_pma_loss_of_signal_o
  , LL_FLOCK_O  => usr_rx1_pma_ll_fast_locked_o
  , LL_SLOCK_O  => usr_rx1_pma_ll_slow_locked_o
  , PLL_LOCK_O  => usr_rx1_pma_pll_lock_o
  , PLL_LOCKT_O => usr_rx1_pma_pll_lock_track_o

  , LINK       => LINK_RX1
);
--#}}}#

-- txlane2: NX_CTX_U#{{{#
txlane2: NX_CTX_U generic map (
   cfg_tx_pcs_protocol_size_i    => cfg_tx2_pcs_protocol_size_i
 , cfg_tx_pcs_8b_scr_sel_i       => cfg_tx2_pcs_8b_scr_sel_i
 , cfg_tx_pcs_scr_init_i         => cfg_tx2_pcs_scr_init_i
 , cfg_tx_pcs_scr_bypass_i       => cfg_tx2_pcs_scr_bypass_i
 , cfg_tx_pcs_sync_supported_i   => cfg_tx2_pcs_sync_supported_i
 , cfg_tx_pcs_replace_bypass_i   => cfg_tx2_pcs_replace_bypass_i
 , cfg_tx_pcs_enc_bypass_i       => cfg_tx2_pcs_enc_bypass_i
 , cfg_tx_pcs_loopback_i         => cfg_tx2_pcs_loopback_i
 , cfg_tx_pcs_polarity_i         => cfg_tx2_pcs_polarity_i
 , cfg_tx_pcs_esistream_fsm_en_i => cfg_tx2_pcs_esistream_fsm_en_i
 , cfg_tx_pcs_bypass_pma_cdc_i   => cfg_tx2_pcs_bypass_pma_cdc_i
 , cfg_tx_pcs_bypass_usr_cdc_i   => cfg_tx2_pcs_bypass_usr_cdc_i
 , cfg_tx_pma_clk_pos_i          => cfg_tx2_pma_clk_pos_i
 , cfg_tx_pma_loopback_i         => cfg_tx2_pma_loopback_i
 , cfg_tx_gearbox_en_i           => cfg_tx2_gearbox_en_i
 , cfg_tx_gearbox_mode_i         => cfg_tx2_gearbox_mode_i
 , location                      => location & ":CHANNEL3.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx2_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx2_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx2_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx2_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx2_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx2_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx2_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx2_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx2_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx2_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx2_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx2_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx2_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx2_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx2_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx2_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx2_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx2_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx2_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx2_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx2_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx2_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx2_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx2_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx2_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx2_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx2_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx2_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx2_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx2_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx2_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx2_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx2_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx2_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx2_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx2_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx2_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx2_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx2_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx2_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx2_ctrl_replace_en_i
  , RST_N_I  => usr_tx2_rst_n_i

  , DATA_I1  => usr_tx2_data_i(0)
  , DATA_I2  => usr_tx2_data_i(1)
  , DATA_I3  => usr_tx2_data_i(2)
  , DATA_I4  => usr_tx2_data_i(3)
  , DATA_I5  => usr_tx2_data_i(4)
  , DATA_I6  => usr_tx2_data_i(5)
  , DATA_I7  => usr_tx2_data_i(6)
  , DATA_I8  => usr_tx2_data_i(7)
  , DATA_I9  => usr_tx2_data_i(8)
  , DATA_I10 => usr_tx2_data_i(9)
  , DATA_I11 => usr_tx2_data_i(10)
  , DATA_I12 => usr_tx2_data_i(11)
  , DATA_I13 => usr_tx2_data_i(12)
  , DATA_I14 => usr_tx2_data_i(13)
  , DATA_I15 => usr_tx2_data_i(14)
  , DATA_I16 => usr_tx2_data_i(15)
  , DATA_I17 => usr_tx2_data_i(16)
  , DATA_I18 => usr_tx2_data_i(17)
  , DATA_I19 => usr_tx2_data_i(18)
  , DATA_I20 => usr_tx2_data_i(19)
  , DATA_I21 => usr_tx2_data_i(20)
  , DATA_I22 => usr_tx2_data_i(21)
  , DATA_I23 => usr_tx2_data_i(22)
  , DATA_I24 => usr_tx2_data_i(23)
  , DATA_I25 => usr_tx2_data_i(24)
  , DATA_I26 => usr_tx2_data_i(25)
  , DATA_I27 => usr_tx2_data_i(26)
  , DATA_I28 => usr_tx2_data_i(27)
  , DATA_I29 => usr_tx2_data_i(28)
  , DATA_I30 => usr_tx2_data_i(29)
  , DATA_I31 => usr_tx2_data_i(30)
  , DATA_I32 => usr_tx2_data_i(31)
  , DATA_I33 => usr_tx2_data_i(32)
  , DATA_I34 => usr_tx2_data_i(33)
  , DATA_I35 => usr_tx2_data_i(34)
  , DATA_I36 => usr_tx2_data_i(35)
  , DATA_I37 => usr_tx2_data_i(36)
  , DATA_I38 => usr_tx2_data_i(37)
  , DATA_I39 => usr_tx2_data_i(38)
  , DATA_I40 => usr_tx2_data_i(39)
  , DATA_I41 => usr_tx2_data_i(40)
  , DATA_I42 => usr_tx2_data_i(41)
  , DATA_I43 => usr_tx2_data_i(42)
  , DATA_I44 => usr_tx2_data_i(43)
  , DATA_I45 => usr_tx2_data_i(44)
  , DATA_I46 => usr_tx2_data_i(45)
  , DATA_I47 => usr_tx2_data_i(46)
  , DATA_I48 => usr_tx2_data_i(47)
  , DATA_I49 => usr_tx2_data_i(48)
  , DATA_I50 => usr_tx2_data_i(49)
  , DATA_I51 => usr_tx2_data_i(50)
  , DATA_I52 => usr_tx2_data_i(51)
  , DATA_I53 => usr_tx2_data_i(52)
  , DATA_I54 => usr_tx2_data_i(53)
  , DATA_I55 => usr_tx2_data_i(54)
  , DATA_I56 => usr_tx2_data_i(55)
  , DATA_I57 => usr_tx2_data_i(56)
  , DATA_I58 => usr_tx2_data_i(57)
  , DATA_I59 => usr_tx2_data_i(58)
  , DATA_I60 => usr_tx2_data_i(59)
  , DATA_I61 => usr_tx2_data_i(60)
  , DATA_I62 => usr_tx2_data_i(61)
  , DATA_I63 => usr_tx2_data_i(62)
  , DATA_I64 => usr_tx2_data_i(63)

  , BUSY_O   => usr_tx2_busy_o
  , INV_K_O  => usr_tx2_ctrl_invalid_k_o

  , PWDN_N_I => usr_tx2_ctrl_driver_pwrdwn_n_i
  , CLK_E_I  => usr_tx2_pma_clk_en_i
  , CLK_O    => usr_tx2_pma_tx_clk_o

  , LINK     => LINK_TX2
);
--#}}}#

-- rxlane2: NX_CRX_U#{{{#
rxlane2: NX_CRX_U generic map (
    cfg_rx_pma_m_eye_ppm_i               => cfg_rx2_pma_m_eye_ppm_i
  , cfg_rx_pma_coarse_ppm_i              => cfg_rx2_pma_coarse_ppm_i
  , cfg_rx_pma_fine_ppm_i                => cfg_rx2_pma_fine_ppm_i
  , cfg_rx_pma_peak_detect_cmd_i         => cfg_rx2_pma_peak_detect_cmd_i
  , cfg_rx_pma_peak_detect_on_i          => cfg_rx2_pma_peak_detect_on_i
  , cfg_rx_pma_dco_reg_res_i             => cfg_rx2_pma_dco_reg_res_i
  , cfg_rx_pma_dco_vref_sel_i            => cfg_rx2_pma_dco_vref_sel_i
  , cfg_rx_pma_dco_divl_i                => cfg_rx2_pma_dco_divl_i
  , cfg_rx_pma_dco_divm_i                => cfg_rx2_pma_dco_divm_i
  , cfg_rx_pma_dco_divn_i                => cfg_rx2_pma_dco_divn_i
  , cfg_rx_pma_loopback_i                => cfg_rx2_pma_loopback_i
  , cfg_rx_pma_clk_pos_i                 => cfg_rx2_pma_clk_pos_i
  , cfg_rx_pma_cdr_cp_i                  => cfg_rx2_pma_cdr_cp_i
  , cfg_rx_pma_ctrl_term_i               => cfg_rx2_pma_ctrl_term_i
  , cfg_rx_pma_pll_divf_en_n_i           => cfg_rx2_pma_pll_divf_en_n_i
  , cfg_rx_pma_pll_divm_en_n_i           => cfg_rx2_pma_pll_divm_en_n_i
  , cfg_rx_pma_pll_divn_en_n_i           => cfg_rx2_pma_pll_divn_en_n_i
  , cfg_rx_pma_pll_cpump_n_i             => cfg_rx2_pma_pll_cpump_n_i
  , cfg_rx_pma_pll_divf_i                => cfg_rx2_pma_pll_divf_i
  , cfg_rx_pma_pll_divm_i                => cfg_rx2_pma_pll_divm_i
  , cfg_rx_pma_pll_divn_i                => cfg_rx2_pma_pll_divn_i
  , cfg_rx_pcs_debug_en_i                => cfg_rx2_pcs_debug_en_i
  , cfg_rx_pcs_bypass_pma_cdc_i          => cfg_rx2_pcs_bypass_pma_cdc_i
  , cfg_rx_pcs_fsm_watchdog_en_i         => cfg_rx2_pcs_fsm_watchdog_en_i
  , cfg_rx_pcs_fsm_sel_i                 => cfg_rx2_pcs_fsm_sel_i
  , cfg_rx_pcs_polarity_i                => cfg_rx2_pcs_polarity_i
  , cfg_rx_pcs_loopback_i                => cfg_rx2_pcs_loopback_i
  , cfg_rx_pcs_dscr_bypass_i             => cfg_rx2_pcs_dscr_bypass_i
  , cfg_rx_pcs_8b_dscr_sel_i             => cfg_rx2_pcs_8b_dscr_sel_i
  , cfg_rx_pcs_replace_bypass_i          => cfg_rx2_pcs_replace_bypass_i
  , cfg_rx_pcs_sync_supported_i          => cfg_rx2_pcs_sync_supported_i
  , cfg_rx_pcs_buffers_bypass_i          => cfg_rx2_pcs_buffers_bypass_i
  , cfg_rx_pcs_buffers_use_cdc_i         => cfg_rx2_pcs_buffers_use_cdc_i
  , cfg_rx_pcs_el_buff_skp_header_3_i    => cfg_rx2_pcs_el_buff_skp_header_3_i
  , cfg_rx_pcs_el_buff_skp_header_2_i    => cfg_rx2_pcs_el_buff_skp_header_2_i
  , cfg_rx_pcs_el_buff_skp_header_1_i    => cfg_rx2_pcs_el_buff_skp_header_1_i
  , cfg_rx_pcs_el_buff_skp_header_0_i    => cfg_rx2_pcs_el_buff_skp_header_0_i
  , cfg_rx_pcs_el_buff_skp_header_size_i => cfg_rx2_pcs_el_buff_skp_header_size_i
  , cfg_rx_pcs_el_buff_skp_char_3_i      => cfg_rx2_pcs_el_buff_skp_char_3_i
  , cfg_rx_pcs_el_buff_skp_char_2_i      => cfg_rx2_pcs_el_buff_skp_char_2_i
  , cfg_rx_pcs_el_buff_skp_char_1_i      => cfg_rx2_pcs_el_buff_skp_char_1_i
  , cfg_rx_pcs_el_buff_skp_char_0_i      => cfg_rx2_pcs_el_buff_skp_char_0_i
  , cfg_rx_pcs_el_buff_skp_seq_size_i    => cfg_rx2_pcs_el_buff_skp_seq_size_i
  , cfg_rx_pcs_el_buff_only_one_skp_i    => cfg_rx2_pcs_el_buff_only_one_skp_i
  , cfg_rx_pcs_el_buff_diff_bef_comp_i   => cfg_rx2_pcs_el_buff_diff_bef_comp_i
  , cfg_rx_pcs_el_buff_max_comp_i        => cfg_rx2_pcs_el_buff_max_comp_i
  , cfg_rx_pcs_dec_bypass_i              => cfg_rx2_pcs_dec_bypass_i
  , cfg_rx_pcs_align_bypass_i            => cfg_rx2_pcs_align_bypass_i
  , cfg_rx_pcs_nb_comma_bef_realign_i    => cfg_rx2_pcs_nb_comma_bef_realign_i
  , cfg_rx_pcs_comma_mask_i              => cfg_rx2_pcs_comma_mask_i
  , cfg_rx_pcs_m_comma_val_i             => cfg_rx2_pcs_m_comma_val_i
  , cfg_rx_pcs_m_comma_en_i              => cfg_rx2_pcs_m_comma_en_i
  , cfg_rx_pcs_p_comma_val_i             => cfg_rx2_pcs_p_comma_val_i
  , cfg_rx_pcs_p_comma_en_i              => cfg_rx2_pcs_p_comma_en_i
  , cfg_rx_pcs_bypass_usr_cdc_i          => cfg_rx2_pcs_bypass_usr_cdc_i
  , cfg_rx_pcs_protocol_size_i           => cfg_rx2_pcs_protocol_size_i
  , cfg_rx_gearbox_mode_i                => cfg_rx2_gearbox_mode_i
  , cfg_rx_gearbox_en_i                  => cfg_rx2_gearbox_en_i
  , location                             => location & ":CHANNEL3.CRX1"
 )
port map (
    DSCR_E_I    => usr_rx2_ctrl_dscr_en_i
  , DEC_E_I     => usr_rx2_ctrl_dec_en_i
  , ALIGN_E_I   => usr_rx2_ctrl_align_en_i
  , ALIGN_S_I   => usr_rx2_ctrl_align_sync_i
  , REP_E_I     => usr_rx2_ctrl_replace_en_i
  , BUF_R_I     => usr_rx2_ctrl_el_buff_rst_i

  , OVS_BS_I1   => usr_rx2_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2   => usr_rx2_ctrl_ovs_bit_sel_i(1)

  , RST_N_I     => usr_rx2_rst_n_i

  , PMA_RSTN_I  => usr_rx2_pma_rst_n_i
  , MEYE_RST_I  => usr_rx2_pma_m_eye_rst_i
  , PWDN_N_I    => usr_rx2_pma_pwr_down_n_i
  , DBG_S_I1    => usr_rx2_ctrl_debug_sel_i(0)
  , DBG_S_I2    => usr_rx2_ctrl_debug_sel_i(1)
  , DBG_S_I3    => usr_rx2_ctrl_debug_sel_i(2)

  , DATA_O1     => usr_rx2_data_o(0)
  , DATA_O2     => usr_rx2_data_o(1)
  , DATA_O3     => usr_rx2_data_o(2)
  , DATA_O4     => usr_rx2_data_o(3)
  , DATA_O5     => usr_rx2_data_o(4)
  , DATA_O6     => usr_rx2_data_o(5)
  , DATA_O7     => usr_rx2_data_o(6)
  , DATA_O8     => usr_rx2_data_o(7)
  , DATA_O9     => usr_rx2_data_o(8)
  , DATA_O10    => usr_rx2_data_o(9)
  , DATA_O11    => usr_rx2_data_o(10)
  , DATA_O12    => usr_rx2_data_o(11)
  , DATA_O13    => usr_rx2_data_o(12)
  , DATA_O14    => usr_rx2_data_o(13)
  , DATA_O15    => usr_rx2_data_o(14)
  , DATA_O16    => usr_rx2_data_o(15)
  , DATA_O17    => usr_rx2_data_o(16)
  , DATA_O18    => usr_rx2_data_o(17)
  , DATA_O19    => usr_rx2_data_o(18)
  , DATA_O20    => usr_rx2_data_o(19)
  , DATA_O21    => usr_rx2_data_o(20)
  , DATA_O22    => usr_rx2_data_o(21)
  , DATA_O23    => usr_rx2_data_o(22)
  , DATA_O24    => usr_rx2_data_o(23)
  , DATA_O25    => usr_rx2_data_o(24)
  , DATA_O26    => usr_rx2_data_o(25)
  , DATA_O27    => usr_rx2_data_o(26)
  , DATA_O28    => usr_rx2_data_o(27)
  , DATA_O29    => usr_rx2_data_o(28)
  , DATA_O30    => usr_rx2_data_o(29)
  , DATA_O31    => usr_rx2_data_o(30)
  , DATA_O32    => usr_rx2_data_o(31)
  , DATA_O33    => usr_rx2_data_o(32)
  , DATA_O34    => usr_rx2_data_o(33)
  , DATA_O35    => usr_rx2_data_o(34)
  , DATA_O36    => usr_rx2_data_o(35)
  , DATA_O37    => usr_rx2_data_o(36)
  , DATA_O38    => usr_rx2_data_o(37)
  , DATA_O39    => usr_rx2_data_o(38)
  , DATA_O40    => usr_rx2_data_o(39)
  , DATA_O41    => usr_rx2_data_o(40)
  , DATA_O42    => usr_rx2_data_o(41)
  , DATA_O43    => usr_rx2_data_o(42)
  , DATA_O44    => usr_rx2_data_o(43)
  , DATA_O45    => usr_rx2_data_o(44)
  , DATA_O46    => usr_rx2_data_o(45)
  , DATA_O47    => usr_rx2_data_o(46)
  , DATA_O48    => usr_rx2_data_o(47)
  , DATA_O49    => usr_rx2_data_o(48)
  , DATA_O50    => usr_rx2_data_o(49)
  , DATA_O51    => usr_rx2_data_o(50)
  , DATA_O52    => usr_rx2_data_o(51)
  , DATA_O53    => usr_rx2_data_o(52)
  , DATA_O54    => usr_rx2_data_o(53)
  , DATA_O55    => usr_rx2_data_o(54)
  , DATA_O56    => usr_rx2_data_o(55)
  , DATA_O57    => usr_rx2_data_o(56)
  , DATA_O58    => usr_rx2_data_o(57)
  , DATA_O59    => usr_rx2_data_o(58)
  , DATA_O60    => usr_rx2_data_o(59)
  , DATA_O61    => usr_rx2_data_o(60)
  , DATA_O62    => usr_rx2_data_o(61)
  , DATA_O63    => usr_rx2_data_o(62)
  , DATA_O64    => usr_rx2_data_o(63)

  , CH_COM_O1   => usr_rx2_ctrl_char_is_comma_o(0)
  , CH_COM_O2   => usr_rx2_ctrl_char_is_comma_o(1)
  , CH_COM_O3   => usr_rx2_ctrl_char_is_comma_o(2)
  , CH_COM_O4   => usr_rx2_ctrl_char_is_comma_o(3)
  , CH_COM_O5   => usr_rx2_ctrl_char_is_comma_o(4)
  , CH_COM_O6   => usr_rx2_ctrl_char_is_comma_o(5)
  , CH_COM_O7   => usr_rx2_ctrl_char_is_comma_o(6)
  , CH_COM_O8   => usr_rx2_ctrl_char_is_comma_o(7)

  , CH_K_O1     => usr_rx2_ctrl_char_is_k_o(0)
  , CH_K_O2     => usr_rx2_ctrl_char_is_k_o(1)
  , CH_K_O3     => usr_rx2_ctrl_char_is_k_o(2)
  , CH_K_O4     => usr_rx2_ctrl_char_is_k_o(3)
  , CH_K_O5     => usr_rx2_ctrl_char_is_k_o(4)
  , CH_K_O6     => usr_rx2_ctrl_char_is_k_o(5)
  , CH_K_O7     => usr_rx2_ctrl_char_is_k_o(6)
  , CH_K_O8     => usr_rx2_ctrl_char_is_k_o(7)

  , NIT_O1      => usr_rx2_ctrl_not_in_table_o(0)
  , NIT_O2      => usr_rx2_ctrl_not_in_table_o(1)
  , NIT_O3      => usr_rx2_ctrl_not_in_table_o(2)
  , NIT_O4      => usr_rx2_ctrl_not_in_table_o(3)
  , NIT_O5      => usr_rx2_ctrl_not_in_table_o(4)
  , NIT_O6      => usr_rx2_ctrl_not_in_table_o(5)
  , NIT_O7      => usr_rx2_ctrl_not_in_table_o(6)
  , NIT_O8      => usr_rx2_ctrl_not_in_table_o(7)

  , D_ERR_O1    => usr_rx2_ctrl_disp_err_o(0)
  , D_ERR_O2    => usr_rx2_ctrl_disp_err_o(1)
  , D_ERR_O3    => usr_rx2_ctrl_disp_err_o(2)
  , D_ERR_O4    => usr_rx2_ctrl_disp_err_o(3)
  , D_ERR_O5    => usr_rx2_ctrl_disp_err_o(4)
  , D_ERR_O6    => usr_rx2_ctrl_disp_err_o(5)
  , D_ERR_O7    => usr_rx2_ctrl_disp_err_o(6)
  , D_ERR_O8    => usr_rx2_ctrl_disp_err_o(7)

  , CH_A_O1     => usr_rx2_ctrl_char_is_a_o(0)
  , CH_A_O2     => usr_rx2_ctrl_char_is_a_o(1)
  , CH_A_O3     => usr_rx2_ctrl_char_is_a_o(2)
  , CH_A_O4     => usr_rx2_ctrl_char_is_a_o(3)
  , CH_A_O5     => usr_rx2_ctrl_char_is_a_o(4)
  , CH_A_O6     => usr_rx2_ctrl_char_is_a_o(5)
  , CH_A_O7     => usr_rx2_ctrl_char_is_a_o(6)
  , CH_A_O8     => usr_rx2_ctrl_char_is_a_o(7)

  , CH_F_O1     => usr_rx2_ctrl_char_is_f_o(0)
  , CH_F_O2     => usr_rx2_ctrl_char_is_f_o(1)
  , CH_F_O3     => usr_rx2_ctrl_char_is_f_o(2)
  , CH_F_O4     => usr_rx2_ctrl_char_is_f_o(3)
  , CH_F_O5     => usr_rx2_ctrl_char_is_f_o(4)
  , CH_F_O6     => usr_rx2_ctrl_char_is_f_o(5)
  , CH_F_O7     => usr_rx2_ctrl_char_is_f_o(6)
  , CH_F_O8     => usr_rx2_ctrl_char_is_f_o(7)

  , ALIGN_O     => usr_rx2_ctrl_char_is_aligned_o
  , VREALIGN_O  => usr_rx2_ctrl_valid_realign_o
  , BUSY_O      => usr_rx2_busy_o

  , TST_O1      => usr_rx2_test_o(0)
  , TST_O2      => usr_rx2_test_o(1)
  , TST_O3      => usr_rx2_test_o(2)
  , TST_O4      => usr_rx2_test_o(3)
  , TST_O5      => usr_rx2_test_o(4)
  , TST_O6      => usr_rx2_test_o(5)
  , TST_O7      => usr_rx2_test_o(6)
  , TST_O8      => usr_rx2_test_o(7)

  , LOS_O       => usr_rx2_pma_loss_of_signal_o
  , LL_FLOCK_O  => usr_rx2_pma_ll_fast_locked_o
  , LL_SLOCK_O  => usr_rx2_pma_ll_slow_locked_o
  , PLL_LOCK_O  => usr_rx2_pma_pll_lock_o
  , PLL_LOCKT_O => usr_rx2_pma_pll_lock_track_o

  , LINK       => LINK_RX2
);
--#}}}#

-- txlane3: NX_CTX_U#{{{#
txlane3: NX_CTX_U generic map (

   cfg_tx_pcs_protocol_size_i    => cfg_tx3_pcs_protocol_size_i
 , cfg_tx_pcs_8b_scr_sel_i       => cfg_tx3_pcs_8b_scr_sel_i
 , cfg_tx_pcs_scr_init_i         => cfg_tx3_pcs_scr_init_i
 , cfg_tx_pcs_scr_bypass_i       => cfg_tx3_pcs_scr_bypass_i
 , cfg_tx_pcs_sync_supported_i   => cfg_tx3_pcs_sync_supported_i
 , cfg_tx_pcs_replace_bypass_i   => cfg_tx3_pcs_replace_bypass_i
 , cfg_tx_pcs_enc_bypass_i       => cfg_tx3_pcs_enc_bypass_i
 , cfg_tx_pcs_loopback_i         => cfg_tx3_pcs_loopback_i
 , cfg_tx_pcs_polarity_i         => cfg_tx3_pcs_polarity_i
 , cfg_tx_pcs_esistream_fsm_en_i => cfg_tx3_pcs_esistream_fsm_en_i
 , cfg_tx_pcs_bypass_pma_cdc_i   => cfg_tx3_pcs_bypass_pma_cdc_i
 , cfg_tx_pcs_bypass_usr_cdc_i   => cfg_tx3_pcs_bypass_usr_cdc_i
 , cfg_tx_pma_clk_pos_i          => cfg_tx3_pma_clk_pos_i
 , cfg_tx_pma_loopback_i         => cfg_tx3_pma_loopback_i
 , cfg_tx_gearbox_en_i           => cfg_tx3_gearbox_en_i
 , cfg_tx_gearbox_mode_i         => cfg_tx3_gearbox_mode_i
 , location                      => location & ":CHANNEL4.CTX1"
 )
port map (
    ENC_E_I1 => usr_tx3_ctrl_enc_en_i(0)
  , ENC_E_I2 => usr_tx3_ctrl_enc_en_i(1)
  , ENC_E_I3 => usr_tx3_ctrl_enc_en_i(2)
  , ENC_E_I4 => usr_tx3_ctrl_enc_en_i(3)
  , ENC_E_I5 => usr_tx3_ctrl_enc_en_i(4)
  , ENC_E_I6 => usr_tx3_ctrl_enc_en_i(5)
  , ENC_E_I7 => usr_tx3_ctrl_enc_en_i(6)
  , ENC_E_I8 => usr_tx3_ctrl_enc_en_i(7)

  , CH_K_I1  => usr_tx3_ctrl_char_is_k_i(0)
  , CH_K_I2  => usr_tx3_ctrl_char_is_k_i(1)
  , CH_K_I3  => usr_tx3_ctrl_char_is_k_i(2)
  , CH_K_I4  => usr_tx3_ctrl_char_is_k_i(3)
  , CH_K_I5  => usr_tx3_ctrl_char_is_k_i(4)
  , CH_K_I6  => usr_tx3_ctrl_char_is_k_i(5)
  , CH_K_I7  => usr_tx3_ctrl_char_is_k_i(6)
  , CH_K_I8  => usr_tx3_ctrl_char_is_k_i(7)

  , SCR_E_I1 => usr_tx3_ctrl_scr_en_i(0)
  , SCR_E_I2 => usr_tx3_ctrl_scr_en_i(1)
  , SCR_E_I3 => usr_tx3_ctrl_scr_en_i(2)
  , SCR_E_I4 => usr_tx3_ctrl_scr_en_i(3)
  , SCR_E_I5 => usr_tx3_ctrl_scr_en_i(4)
  , SCR_E_I6 => usr_tx3_ctrl_scr_en_i(5)
  , SCR_E_I7 => usr_tx3_ctrl_scr_en_i(6)
  , SCR_E_I8 => usr_tx3_ctrl_scr_en_i(7)

  , EOMF_I1  => usr_tx3_ctrl_end_of_multiframe_i(0)
  , EOMF_I2  => usr_tx3_ctrl_end_of_multiframe_i(1)
  , EOMF_I3  => usr_tx3_ctrl_end_of_multiframe_i(2)
  , EOMF_I4  => usr_tx3_ctrl_end_of_multiframe_i(3)
  , EOMF_I5  => usr_tx3_ctrl_end_of_multiframe_i(4)
  , EOMF_I6  => usr_tx3_ctrl_end_of_multiframe_i(5)
  , EOMF_I7  => usr_tx3_ctrl_end_of_multiframe_i(6)
  , EOMF_I8  => usr_tx3_ctrl_end_of_multiframe_i(7)

  , EOF_I1   => usr_tx3_ctrl_end_of_frame_i(0)
  , EOF_I2   => usr_tx3_ctrl_end_of_frame_i(1)
  , EOF_I3   => usr_tx3_ctrl_end_of_frame_i(2)
  , EOF_I4   => usr_tx3_ctrl_end_of_frame_i(3)
  , EOF_I5   => usr_tx3_ctrl_end_of_frame_i(4)
  , EOF_I6   => usr_tx3_ctrl_end_of_frame_i(5)
  , EOF_I7   => usr_tx3_ctrl_end_of_frame_i(6)
  , EOF_I8   => usr_tx3_ctrl_end_of_frame_i(7)

  , REP_E_I  => usr_tx3_ctrl_replace_en_i
  , RST_N_I  => usr_tx3_rst_n_i

  , DATA_I1  => usr_tx3_data_i(0)
  , DATA_I2  => usr_tx3_data_i(1)
  , DATA_I3  => usr_tx3_data_i(2)
  , DATA_I4  => usr_tx3_data_i(3)
  , DATA_I5  => usr_tx3_data_i(4)
  , DATA_I6  => usr_tx3_data_i(5)
  , DATA_I7  => usr_tx3_data_i(6)
  , DATA_I8  => usr_tx3_data_i(7)
  , DATA_I9  => usr_tx3_data_i(8)
  , DATA_I10 => usr_tx3_data_i(9)
  , DATA_I11 => usr_tx3_data_i(10)
  , DATA_I12 => usr_tx3_data_i(11)
  , DATA_I13 => usr_tx3_data_i(12)
  , DATA_I14 => usr_tx3_data_i(13)
  , DATA_I15 => usr_tx3_data_i(14)
  , DATA_I16 => usr_tx3_data_i(15)
  , DATA_I17 => usr_tx3_data_i(16)
  , DATA_I18 => usr_tx3_data_i(17)
  , DATA_I19 => usr_tx3_data_i(18)
  , DATA_I20 => usr_tx3_data_i(19)
  , DATA_I21 => usr_tx3_data_i(20)
  , DATA_I22 => usr_tx3_data_i(21)
  , DATA_I23 => usr_tx3_data_i(22)
  , DATA_I24 => usr_tx3_data_i(23)
  , DATA_I25 => usr_tx3_data_i(24)
  , DATA_I26 => usr_tx3_data_i(25)
  , DATA_I27 => usr_tx3_data_i(26)
  , DATA_I28 => usr_tx3_data_i(27)
  , DATA_I29 => usr_tx3_data_i(28)
  , DATA_I30 => usr_tx3_data_i(29)
  , DATA_I31 => usr_tx3_data_i(30)
  , DATA_I32 => usr_tx3_data_i(31)
  , DATA_I33 => usr_tx3_data_i(32)
  , DATA_I34 => usr_tx3_data_i(33)
  , DATA_I35 => usr_tx3_data_i(34)
  , DATA_I36 => usr_tx3_data_i(35)
  , DATA_I37 => usr_tx3_data_i(36)
  , DATA_I38 => usr_tx3_data_i(37)
  , DATA_I39 => usr_tx3_data_i(38)
  , DATA_I40 => usr_tx3_data_i(39)
  , DATA_I41 => usr_tx3_data_i(40)
  , DATA_I42 => usr_tx3_data_i(41)
  , DATA_I43 => usr_tx3_data_i(42)
  , DATA_I44 => usr_tx3_data_i(43)
  , DATA_I45 => usr_tx3_data_i(44)
  , DATA_I46 => usr_tx3_data_i(45)
  , DATA_I47 => usr_tx3_data_i(46)
  , DATA_I48 => usr_tx3_data_i(47)
  , DATA_I49 => usr_tx3_data_i(48)
  , DATA_I50 => usr_tx3_data_i(49)
  , DATA_I51 => usr_tx3_data_i(50)
  , DATA_I52 => usr_tx3_data_i(51)
  , DATA_I53 => usr_tx3_data_i(52)
  , DATA_I54 => usr_tx3_data_i(53)
  , DATA_I55 => usr_tx3_data_i(54)
  , DATA_I56 => usr_tx3_data_i(55)
  , DATA_I57 => usr_tx3_data_i(56)
  , DATA_I58 => usr_tx3_data_i(57)
  , DATA_I59 => usr_tx3_data_i(58)
  , DATA_I60 => usr_tx3_data_i(59)
  , DATA_I61 => usr_tx3_data_i(60)
  , DATA_I62 => usr_tx3_data_i(61)
  , DATA_I63 => usr_tx3_data_i(62)
  , DATA_I64 => usr_tx3_data_i(63)

  , BUSY_O   => usr_tx3_busy_o
  , INV_K_O  => usr_tx3_ctrl_invalid_k_o

  , PWDN_N_I => usr_tx3_ctrl_driver_pwrdwn_n_i
  , CLK_E_I  => usr_tx3_pma_clk_en_i
  , CLK_O    => usr_tx3_pma_tx_clk_o

  , LINK     => LINK_TX3
);
--#}}}#

-- rxlane3: NX_CRX_U#{{{#
rxlane3: NX_CRX_U generic map (
    cfg_rx_pma_m_eye_ppm_i               => cfg_rx3_pma_m_eye_ppm_i
  , cfg_rx_pma_coarse_ppm_i              => cfg_rx3_pma_coarse_ppm_i
  , cfg_rx_pma_fine_ppm_i                => cfg_rx3_pma_fine_ppm_i
  , cfg_rx_pma_peak_detect_cmd_i         => cfg_rx3_pma_peak_detect_cmd_i
  , cfg_rx_pma_peak_detect_on_i          => cfg_rx3_pma_peak_detect_on_i
  , cfg_rx_pma_dco_reg_res_i             => cfg_rx3_pma_dco_reg_res_i
  , cfg_rx_pma_dco_vref_sel_i            => cfg_rx3_pma_dco_vref_sel_i
  , cfg_rx_pma_dco_divl_i                => cfg_rx3_pma_dco_divl_i
  , cfg_rx_pma_dco_divm_i                => cfg_rx3_pma_dco_divm_i
  , cfg_rx_pma_dco_divn_i                => cfg_rx3_pma_dco_divn_i
  , cfg_rx_pma_loopback_i                => cfg_rx3_pma_loopback_i
  , cfg_rx_pma_clk_pos_i                 => cfg_rx3_pma_clk_pos_i
  , cfg_rx_pma_cdr_cp_i                  => cfg_rx3_pma_cdr_cp_i
  , cfg_rx_pma_ctrl_term_i               => cfg_rx3_pma_ctrl_term_i
  , cfg_rx_pma_pll_divf_en_n_i           => cfg_rx3_pma_pll_divf_en_n_i
  , cfg_rx_pma_pll_divm_en_n_i           => cfg_rx3_pma_pll_divm_en_n_i
  , cfg_rx_pma_pll_divn_en_n_i           => cfg_rx3_pma_pll_divn_en_n_i
  , cfg_rx_pma_pll_cpump_n_i             => cfg_rx3_pma_pll_cpump_n_i
  , cfg_rx_pma_pll_divf_i                => cfg_rx3_pma_pll_divf_i
  , cfg_rx_pma_pll_divm_i                => cfg_rx3_pma_pll_divm_i
  , cfg_rx_pma_pll_divn_i                => cfg_rx3_pma_pll_divn_i
  , cfg_rx_pcs_debug_en_i                => cfg_rx3_pcs_debug_en_i
  , cfg_rx_pcs_bypass_pma_cdc_i          => cfg_rx3_pcs_bypass_pma_cdc_i
  , cfg_rx_pcs_fsm_watchdog_en_i         => cfg_rx3_pcs_fsm_watchdog_en_i
  , cfg_rx_pcs_fsm_sel_i                 => cfg_rx3_pcs_fsm_sel_i
  , cfg_rx_pcs_polarity_i                => cfg_rx3_pcs_polarity_i
  , cfg_rx_pcs_loopback_i                => cfg_rx3_pcs_loopback_i
  , cfg_rx_pcs_dscr_bypass_i             => cfg_rx3_pcs_dscr_bypass_i
  , cfg_rx_pcs_8b_dscr_sel_i             => cfg_rx3_pcs_8b_dscr_sel_i
  , cfg_rx_pcs_replace_bypass_i          => cfg_rx3_pcs_replace_bypass_i
  , cfg_rx_pcs_sync_supported_i          => cfg_rx3_pcs_sync_supported_i
  , cfg_rx_pcs_buffers_bypass_i          => cfg_rx3_pcs_buffers_bypass_i
  , cfg_rx_pcs_buffers_use_cdc_i         => cfg_rx3_pcs_buffers_use_cdc_i
  , cfg_rx_pcs_el_buff_skp_header_3_i    => cfg_rx3_pcs_el_buff_skp_header_3_i
  , cfg_rx_pcs_el_buff_skp_header_2_i    => cfg_rx3_pcs_el_buff_skp_header_2_i
  , cfg_rx_pcs_el_buff_skp_header_1_i    => cfg_rx3_pcs_el_buff_skp_header_1_i
  , cfg_rx_pcs_el_buff_skp_header_0_i    => cfg_rx3_pcs_el_buff_skp_header_0_i
  , cfg_rx_pcs_el_buff_skp_header_size_i => cfg_rx3_pcs_el_buff_skp_header_size_i
  , cfg_rx_pcs_el_buff_skp_char_3_i      => cfg_rx3_pcs_el_buff_skp_char_3_i
  , cfg_rx_pcs_el_buff_skp_char_2_i      => cfg_rx3_pcs_el_buff_skp_char_2_i
  , cfg_rx_pcs_el_buff_skp_char_1_i      => cfg_rx3_pcs_el_buff_skp_char_1_i
  , cfg_rx_pcs_el_buff_skp_char_0_i      => cfg_rx3_pcs_el_buff_skp_char_0_i
  , cfg_rx_pcs_el_buff_skp_seq_size_i    => cfg_rx3_pcs_el_buff_skp_seq_size_i
  , cfg_rx_pcs_el_buff_only_one_skp_i    => cfg_rx3_pcs_el_buff_only_one_skp_i
  , cfg_rx_pcs_el_buff_diff_bef_comp_i   => cfg_rx3_pcs_el_buff_diff_bef_comp_i
  , cfg_rx_pcs_el_buff_max_comp_i        => cfg_rx3_pcs_el_buff_max_comp_i
  , cfg_rx_pcs_dec_bypass_i              => cfg_rx3_pcs_dec_bypass_i
  , cfg_rx_pcs_align_bypass_i            => cfg_rx3_pcs_align_bypass_i
  , cfg_rx_pcs_nb_comma_bef_realign_i    => cfg_rx3_pcs_nb_comma_bef_realign_i
  , cfg_rx_pcs_comma_mask_i              => cfg_rx3_pcs_comma_mask_i
  , cfg_rx_pcs_m_comma_val_i             => cfg_rx3_pcs_m_comma_val_i
  , cfg_rx_pcs_m_comma_en_i              => cfg_rx3_pcs_m_comma_en_i
  , cfg_rx_pcs_p_comma_val_i             => cfg_rx3_pcs_p_comma_val_i
  , cfg_rx_pcs_p_comma_en_i              => cfg_rx3_pcs_p_comma_en_i
  , cfg_rx_pcs_bypass_usr_cdc_i          => cfg_rx3_pcs_bypass_usr_cdc_i
  , cfg_rx_pcs_protocol_size_i           => cfg_rx3_pcs_protocol_size_i
  , cfg_rx_gearbox_mode_i                => cfg_rx3_gearbox_mode_i
  , cfg_rx_gearbox_en_i                  => cfg_rx3_gearbox_en_i
  , location                             => location & ":CHANNEL4.CRX1"
 )
port map (
    DSCR_E_I    => usr_rx3_ctrl_dscr_en_i
  , DEC_E_I     => usr_rx3_ctrl_dec_en_i
  , ALIGN_E_I   => usr_rx3_ctrl_align_en_i
  , ALIGN_S_I   => usr_rx3_ctrl_align_sync_i
  , REP_E_I     => usr_rx3_ctrl_replace_en_i
  , BUF_R_I     => usr_rx3_ctrl_el_buff_rst_i

  , OVS_BS_I1   => usr_rx3_ctrl_ovs_bit_sel_i(0)
  , OVS_BS_I2   => usr_rx3_ctrl_ovs_bit_sel_i(1)

  , RST_N_I     => usr_rx3_rst_n_i

  , PMA_RSTN_I  => usr_rx3_pma_rst_n_i
  , MEYE_RST_I  => usr_rx3_pma_m_eye_rst_i
  , PWDN_N_I    => usr_rx3_pma_pwr_down_n_i
  , DBG_S_I1    => usr_rx3_ctrl_debug_sel_i(0)
  , DBG_S_I2    => usr_rx3_ctrl_debug_sel_i(1)
  , DBG_S_I3    => usr_rx3_ctrl_debug_sel_i(2)

  , DATA_O1     => usr_rx3_data_o(0)
  , DATA_O2     => usr_rx3_data_o(1)
  , DATA_O3     => usr_rx3_data_o(2)
  , DATA_O4     => usr_rx3_data_o(3)
  , DATA_O5     => usr_rx3_data_o(4)
  , DATA_O6     => usr_rx3_data_o(5)
  , DATA_O7     => usr_rx3_data_o(6)
  , DATA_O8     => usr_rx3_data_o(7)
  , DATA_O9     => usr_rx3_data_o(8)
  , DATA_O10    => usr_rx3_data_o(9)
  , DATA_O11    => usr_rx3_data_o(10)
  , DATA_O12    => usr_rx3_data_o(11)
  , DATA_O13    => usr_rx3_data_o(12)
  , DATA_O14    => usr_rx3_data_o(13)
  , DATA_O15    => usr_rx3_data_o(14)
  , DATA_O16    => usr_rx3_data_o(15)
  , DATA_O17    => usr_rx3_data_o(16)
  , DATA_O18    => usr_rx3_data_o(17)
  , DATA_O19    => usr_rx3_data_o(18)
  , DATA_O20    => usr_rx3_data_o(19)
  , DATA_O21    => usr_rx3_data_o(20)
  , DATA_O22    => usr_rx3_data_o(21)
  , DATA_O23    => usr_rx3_data_o(22)
  , DATA_O24    => usr_rx3_data_o(23)
  , DATA_O25    => usr_rx3_data_o(24)
  , DATA_O26    => usr_rx3_data_o(25)
  , DATA_O27    => usr_rx3_data_o(26)
  , DATA_O28    => usr_rx3_data_o(27)
  , DATA_O29    => usr_rx3_data_o(28)
  , DATA_O30    => usr_rx3_data_o(29)
  , DATA_O31    => usr_rx3_data_o(30)
  , DATA_O32    => usr_rx3_data_o(31)
  , DATA_O33    => usr_rx3_data_o(32)
  , DATA_O34    => usr_rx3_data_o(33)
  , DATA_O35    => usr_rx3_data_o(34)
  , DATA_O36    => usr_rx3_data_o(35)
  , DATA_O37    => usr_rx3_data_o(36)
  , DATA_O38    => usr_rx3_data_o(37)
  , DATA_O39    => usr_rx3_data_o(38)
  , DATA_O40    => usr_rx3_data_o(39)
  , DATA_O41    => usr_rx3_data_o(40)
  , DATA_O42    => usr_rx3_data_o(41)
  , DATA_O43    => usr_rx3_data_o(42)
  , DATA_O44    => usr_rx3_data_o(43)
  , DATA_O45    => usr_rx3_data_o(44)
  , DATA_O46    => usr_rx3_data_o(45)
  , DATA_O47    => usr_rx3_data_o(46)
  , DATA_O48    => usr_rx3_data_o(47)
  , DATA_O49    => usr_rx3_data_o(48)
  , DATA_O50    => usr_rx3_data_o(49)
  , DATA_O51    => usr_rx3_data_o(50)
  , DATA_O52    => usr_rx3_data_o(51)
  , DATA_O53    => usr_rx3_data_o(52)
  , DATA_O54    => usr_rx3_data_o(53)
  , DATA_O55    => usr_rx3_data_o(54)
  , DATA_O56    => usr_rx3_data_o(55)
  , DATA_O57    => usr_rx3_data_o(56)
  , DATA_O58    => usr_rx3_data_o(57)
  , DATA_O59    => usr_rx3_data_o(58)
  , DATA_O60    => usr_rx3_data_o(59)
  , DATA_O61    => usr_rx3_data_o(60)
  , DATA_O62    => usr_rx3_data_o(61)
  , DATA_O63    => usr_rx3_data_o(62)
  , DATA_O64    => usr_rx3_data_o(63)

  , CH_COM_O1   => usr_rx3_ctrl_char_is_comma_o(0)
  , CH_COM_O2   => usr_rx3_ctrl_char_is_comma_o(1)
  , CH_COM_O3   => usr_rx3_ctrl_char_is_comma_o(2)
  , CH_COM_O4   => usr_rx3_ctrl_char_is_comma_o(3)
  , CH_COM_O5   => usr_rx3_ctrl_char_is_comma_o(4)
  , CH_COM_O6   => usr_rx3_ctrl_char_is_comma_o(5)
  , CH_COM_O7   => usr_rx3_ctrl_char_is_comma_o(6)
  , CH_COM_O8   => usr_rx3_ctrl_char_is_comma_o(7)

  , CH_K_O1     => usr_rx3_ctrl_char_is_k_o(0)
  , CH_K_O2     => usr_rx3_ctrl_char_is_k_o(1)
  , CH_K_O3     => usr_rx3_ctrl_char_is_k_o(2)
  , CH_K_O4     => usr_rx3_ctrl_char_is_k_o(3)
  , CH_K_O5     => usr_rx3_ctrl_char_is_k_o(4)
  , CH_K_O6     => usr_rx3_ctrl_char_is_k_o(5)
  , CH_K_O7     => usr_rx3_ctrl_char_is_k_o(6)
  , CH_K_O8     => usr_rx3_ctrl_char_is_k_o(7)

  , NIT_O1      => usr_rx3_ctrl_not_in_table_o(0)
  , NIT_O2      => usr_rx3_ctrl_not_in_table_o(1)
  , NIT_O3      => usr_rx3_ctrl_not_in_table_o(2)
  , NIT_O4      => usr_rx3_ctrl_not_in_table_o(3)
  , NIT_O5      => usr_rx3_ctrl_not_in_table_o(4)
  , NIT_O6      => usr_rx3_ctrl_not_in_table_o(5)
  , NIT_O7      => usr_rx3_ctrl_not_in_table_o(6)
  , NIT_O8      => usr_rx3_ctrl_not_in_table_o(7)

  , D_ERR_O1    => usr_rx3_ctrl_disp_err_o(0)
  , D_ERR_O2    => usr_rx3_ctrl_disp_err_o(1)
  , D_ERR_O3    => usr_rx3_ctrl_disp_err_o(2)
  , D_ERR_O4    => usr_rx3_ctrl_disp_err_o(3)
  , D_ERR_O5    => usr_rx3_ctrl_disp_err_o(4)
  , D_ERR_O6    => usr_rx3_ctrl_disp_err_o(5)
  , D_ERR_O7    => usr_rx3_ctrl_disp_err_o(6)
  , D_ERR_O8    => usr_rx3_ctrl_disp_err_o(7)

  , CH_A_O1     => usr_rx3_ctrl_char_is_a_o(0)
  , CH_A_O2     => usr_rx3_ctrl_char_is_a_o(1)
  , CH_A_O3     => usr_rx3_ctrl_char_is_a_o(2)
  , CH_A_O4     => usr_rx3_ctrl_char_is_a_o(3)
  , CH_A_O5     => usr_rx3_ctrl_char_is_a_o(4)
  , CH_A_O6     => usr_rx3_ctrl_char_is_a_o(5)
  , CH_A_O7     => usr_rx3_ctrl_char_is_a_o(6)
  , CH_A_O8     => usr_rx3_ctrl_char_is_a_o(7)

  , CH_F_O1     => usr_rx3_ctrl_char_is_f_o(0)
  , CH_F_O2     => usr_rx3_ctrl_char_is_f_o(1)
  , CH_F_O3     => usr_rx3_ctrl_char_is_f_o(2)
  , CH_F_O4     => usr_rx3_ctrl_char_is_f_o(3)
  , CH_F_O5     => usr_rx3_ctrl_char_is_f_o(4)
  , CH_F_O6     => usr_rx3_ctrl_char_is_f_o(5)
  , CH_F_O7     => usr_rx3_ctrl_char_is_f_o(6)
  , CH_F_O8     => usr_rx3_ctrl_char_is_f_o(7)

  , ALIGN_O     => usr_rx3_ctrl_char_is_aligned_o
  , VREALIGN_O  => usr_rx3_ctrl_valid_realign_o
  , BUSY_O      => usr_rx3_busy_o

  , TST_O1      => usr_rx3_test_o(0)
  , TST_O2      => usr_rx3_test_o(1)
  , TST_O3      => usr_rx3_test_o(2)
  , TST_O4      => usr_rx3_test_o(3)
  , TST_O5      => usr_rx3_test_o(4)
  , TST_O6      => usr_rx3_test_o(5)
  , TST_O7      => usr_rx3_test_o(6)
  , TST_O8      => usr_rx3_test_o(7)

  , LOS_O       => usr_rx3_pma_loss_of_signal_o
  , LL_FLOCK_O  => usr_rx3_pma_ll_fast_locked_o
  , LL_SLOCK_O  => usr_rx3_pma_ll_slow_locked_o
  , PLL_LOCK_O  => usr_rx3_pma_pll_lock_o
  , PLL_LOCKT_O => usr_rx3_pma_pll_lock_track_o

  , LINK       => LINK_RX3
);
--#}}}#

end NX_RTL;
--#}}}#
-- =================================================================================================
--   NX_PMA_U definition                                                                2018/11/30
-- =================================================================================================

-- NX_PMA_U#{{{#
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_PMA_U is
 generic (
   cfg_pll_pma_int_data_len_i            : bit := '0';
   cfg_pll_pma_cpump_i                   : bit_vector( 3 downto 0) := (others => '0');
   cfg_pll_pma_divl_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_divm_i                    : bit := '0';
   cfg_pll_pma_divn_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pll_pma_lvds_en_i                 : bit := '0';
   cfg_pll_pma_lvds_mux_i                : bit := '0';
   cfg_pll_pma_mux_ckref_i               : bit := '0';
   cfg_pll_pma_gbx_en_i                  : bit := '0';
   cfg_pll_pma_ckref_ext_i               : bit := '0';
   cfg_main_clk_to_fabric_div_mode_i     : bit := '0';
   cfg_main_clk_to_fabric_div_en_i       : bit := '0';
   cfg_main_clk_to_fabric_sel_i          : bit := '0';
   cfg_main_rclk_to_fabric_sel_i         : bit_vector( 1 downto 0) := (others => '0');
   cfg_main_use_only_usr_clock_i         : bit := '0';
   tx_usrclk_use_pcs_clk_2               : bit := '0';
   rx_usrclk_use_pcs_clk_2               : bit := '0';
   cfg_pcs_word_len_i                    : bit_vector( 1 downto 0) := (others => '0');
   cfg_pcs_ovs_en_i                      : bit := '0';
   cfg_pcs_ovs_mode_i                    : bit := '0';
   cfg_pcs_pll_lock_ppm_i                : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_m_eye_i            : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_up_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_dn_i         : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_coarse_ena_i : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_fine_ena_i   : bit := '0';
   cfg_dyn_all_rx_pma_m_eye_step_i       : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_mode_i        : bit_vector( 1 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_locked_i      : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_trim_unlocked_i    : bit_vector( 2 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_1        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_all_rx_pma_threshold_2        : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx1_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx2_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx3_pma_pre_sign_i            : bit := '0';
   cfg_dyn_tx0_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx1_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx2_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx3_pma_pre_en_i              : bit := '0';
   cfg_dyn_tx0_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_pre_sel_i             : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_main_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_main_en_i             : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_sel_i          : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_margin_input_i        : bit_vector( 8 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx1_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx2_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx3_pma_post_sign_i           : bit := '0';
   cfg_dyn_tx0_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_en_i             : bit_vector( 4 downto 0) := (others => '0');
   cfg_dyn_tx0_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx1_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx2_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_tx3_pma_post_sel_i            : bit_vector( 7 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_cap_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_ctle_res_p_i          : bit_vector( 3 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap1_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap2_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap3_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_dfe_idac_tap4_n_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx0_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx1_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx2_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_dyn_rx3_pma_termination_cmd_i     : bit_vector( 5 downto 0) := (others => '0');
   cfg_test_mode_i                       : bit_vector( 1 downto 0) := (others => '0');

   location                    : string := ""
);
port (
    CLK_TX_I    : in  std_logic;
    CLK_RX_I    : in  std_logic;
    CLK_REF_I   : in  std_logic;

    DC_E_I       : in  std_logic;
    DC_LCSN_I1   : in  std_logic;
    DC_LCSN_I2   : in  std_logic;
    DC_LCSN_I3   : in  std_logic;
    DC_LCSN_I4   : in  std_logic;

    DC_CCSN_I    : in  std_logic;
    DC_WE_N_I    : in  std_logic;

    DC_ADD_I1    : in  std_logic;
    DC_ADD_I2    : in  std_logic;
    DC_ADD_I3    : in  std_logic;
    DC_ADD_I4    : in  std_logic;
    DC_WDATAS_I  : in  std_logic;
    DC_WDATA_I1  : in  std_logic;
    DC_WDATA_I2  : in  std_logic;
    DC_WDATA_I3  : in  std_logic;
    DC_WDATA_I4  : in  std_logic;
    DC_WDATA_I5  : in  std_logic;
    DC_WDATA_I6  : in  std_logic;
    DC_WDATA_I7  : in  std_logic;
    DC_WDATA_I8  : in  std_logic;
    DC_WDATA_I9  : in  std_logic;
    DC_WDATA_I10 : in  std_logic;
    DC_WDATA_I11 : in  std_logic;
    DC_WDATA_I12 : in  std_logic;

    PLL_RN_I     : in  std_logic;
    PWDN_N_I     : in  std_logic;
    RST_N_I      : in  std_logic;

    DBG_S_I1     : in  std_logic;
    DBG_S_I2     : in  std_logic;
    DBG_A_I      : in  std_logic;

    SE_I         : in  std_logic;

    SCAN_I1      : in  std_logic;
    SCAN_I2      : in  std_logic;
    SCAN_I3      : in  std_logic;
    SCAN_I4      : in  std_logic;
    SCAN_I5      : in  std_logic;
    SCAN_I6      : in  std_logic;
    SCAN_I7      : in  std_logic;
    SCAN_I8      : in  std_logic;

    CLK_O       : out std_logic;
    CLK_RX_O    : out std_logic;
    LOCK_O      : out std_logic;
    LOCKA_O     : out std_logic;
    FB_LOCK_O   : out std_logic;
    CAL_OUT_O   : out std_logic;
    DBG_R_O     : out std_logic;

    LL_O1       : out std_logic;
    LL_O2       : out std_logic;
    LL_O3       : out std_logic;
    LL_O4       : out std_logic;
    LL_O5       : out std_logic;
    LL_O6       : out std_logic;
    LL_O7       : out std_logic;
    LL_O8       : out std_logic;
    LL_O9       : out std_logic;
    LL_O10      : out std_logic;
    LL_O11      : out std_logic;
    LL_O12      : out std_logic;
    LL_O13      : out std_logic;
    LL_O14      : out std_logic;
    LL_O15      : out std_logic;
    LL_O16      : out std_logic;
    LL_O17      : out std_logic;
    LL_O18      : out std_logic;
    LL_O19      : out std_logic;
    LL_O20      : out std_logic;


    SCAN_O1     : out std_logic;
    SCAN_O2     : out std_logic;
    SCAN_O3     : out std_logic;
    SCAN_O4     : out std_logic;
    SCAN_O5     : out std_logic;
    SCAN_O6     : out std_logic;
    SCAN_O7     : out std_logic;
    SCAN_O8     : out std_logic;


    LINK_TX0    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX1    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX2    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_TX3    : inout std_logic_vector(CTX_LINK_SIZE-1 downto 0);
    LINK_RX0    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX1    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX2    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0);
    LINK_RX3    : inout std_logic_vector(CRX_LINK_SIZE-1 downto 0)
);
end NX_PMA_U;
--#}}}#
-- =================================================================================================
--   NX_IOM_L definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_L is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk1 : bit := '0';
--  latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk2 : bit := '0';
--  latency2     : bit := '0';
--  sel_clk_out2 : bit_vector(1 downto 0) := "00";
--  sel_clk_out3 : bit_vector(1 downto 0) := "00";
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_io_cal  : bit := '0';
    pads_dict    : string := "";
    pads_path    : string := ""
);
port(
    RTCK1   : in    std_logic;
    RRCK1   : in    std_logic;
    WTCK1   : in    std_logic;
    WRCK1   : in    std_logic;
    RTCK2   : in    std_logic;
    RRCK2   : in    std_logic;
    WTCK2   : in    std_logic;
    WRCK2   : in    std_logic;
    CTCK    : in    std_logic;
    CCK     : in    std_logic;
    DCK     : in    std_logic;

    C1TW    : in    std_logic;
    C1TS    : in    std_logic;
    C1RW1   : in    std_logic;
    C1RW2   : in    std_logic;
    C1RW3   : in    std_logic;
    C1RNE   : in    std_logic;
    C1RS    : in    std_logic;
    C2TW    : in    std_logic;
    C2TS    : in    std_logic;
    C2RW1   : in    std_logic;
    C2RW2   : in    std_logic;
    C2RW3   : in    std_logic;
    C2RNE   : in    std_logic;
    C2RS    : in    std_logic;
    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;
    DC      : in    std_logic;
    DRI1    : in    std_logic;
    DRI2    : in    std_logic;
    DRI3    : in    std_logic;
    DRI4    : in    std_logic;
    DRI5    : in    std_logic;
    DRI6    : in    std_logic;
    DRA1    : in    std_logic;
    DRA2    : in    std_logic;
    DRA3    : in    std_logic;
    DRA4    : in    std_logic;
    DRA5    : in    std_logic;
    DRA6    : in    std_logic;
    DRL     : in    std_logic;
    DOS     : in    std_logic;
    DOG     : in    std_logic;
    DIS     : in    std_logic;
    DIG     : in    std_logic;
    DPAS    : in    std_logic;
    DPAG    : in    std_logic;
    DQSS    : in    std_logic;
    DQSG    : in    std_logic;
    DS1     : in    std_logic;
    DS2     : in    std_logic;
    CAD1    : in    std_logic;
    CAD2    : in    std_logic;
    CAD3    : in    std_logic;
    CAD4    : in    std_logic;
    CAD5    : in    std_logic;
    CAD6    : in    std_logic;
    CAP1    : in    std_logic;
    CAP2    : in    std_logic;
    CAP3    : in    std_logic;
    CAP4    : in    std_logic;
    CAN1    : in    std_logic;
    CAN2    : in    std_logic;
    CAN3    : in    std_logic;
    CAN4    : in    std_logic;
    CAT1    : in    std_logic;
    CAT2    : in    std_logic;
    CAT3    : in    std_logic;
    CAT4    : in    std_logic;

    CKO1    : out   std_logic;
    CKO2    : out   std_logic;

    FLD     : out   std_logic;
    FLG     : out   std_logic;
    C1RED   : out   std_logic;
    C2RED   : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;
    CAL     : out   std_logic;

    P1CI1   : in    std_logic;
    P1CL    : in    std_logic;
    P1CR    : in    std_logic;
    P1CO    : out   std_logic;
    P1CTI   : in    std_logic;
    P1CTO   : out   std_logic;
    P1EI1   : in    std_logic;
    P1EI2   : in    std_logic;
    P1EI3   : in    std_logic;
    P1EI4   : in    std_logic;
    P1EI5   : in    std_logic;
    P1EL    : in    std_logic;
    P1ER    : in    std_logic;
    P1EO    : out   std_logic;
    P1RI    : in    std_logic;
    P1RL    : in    std_logic;
    P1RR    : in    std_logic;
    P1RO1   : out   std_logic;
    P1RO2   : out   std_logic;
    P1RO3   : out   std_logic;
    P1RO4   : out   std_logic;
    P1RO5   : out   std_logic;

    P2CI1   : in    std_logic;
    P2CL    : in    std_logic;
    P2CR    : in    std_logic;
    P2CO    : out   std_logic;
    P2CTI   : in    std_logic;
    P2CTO   : out   std_logic;
    P2EI1   : in    std_logic;
    P2EI2   : in    std_logic;
    P2EI3   : in    std_logic;
    P2EI4   : in    std_logic;
    P2EI5   : in    std_logic;
    P2EL    : in    std_logic;
    P2ER    : in    std_logic;
    P2EO    : out   std_logic;
    P2RI    : in    std_logic;
    P2RL    : in    std_logic;
    P2RR    : in    std_logic;
    P2RO1   : out   std_logic;
    P2RO2   : out   std_logic;
    P2RO3   : out   std_logic;
    P2RO4   : out   std_logic;
    P2RO5   : out   std_logic;

    P3CI1   : in    std_logic;
    P3CL    : in    std_logic;
    P3CR    : in    std_logic;
    P3CO    : out   std_logic;
    P3CTI   : in    std_logic;
    P3CTO   : out   std_logic;
    P3EI1   : in    std_logic;
    P3EI2   : in    std_logic;
    P3EI3   : in    std_logic;
    P3EI4   : in    std_logic;
    P3EI5   : in    std_logic;
    P3EL    : in    std_logic;
    P3ER    : in    std_logic;
    P3EO    : out   std_logic;
    P3RI    : in    std_logic;
    P3RL    : in    std_logic;
    P3RR    : in    std_logic;
    P3RO1   : out   std_logic;
    P3RO2   : out   std_logic;
    P3RO3   : out   std_logic;
    P3RO4   : out   std_logic;
    P3RO5   : out   std_logic;

    P4CI1   : in    std_logic;
    P4CL    : in    std_logic;
    P4CR    : in    std_logic;
    P4CO    : out   std_logic;
    P4CTI   : in    std_logic;
    P4CTO   : out   std_logic;
    P4EI1   : in    std_logic;
    P4EI2   : in    std_logic;
    P4EI3   : in    std_logic;
    P4EI4   : in    std_logic;
    P4EI5   : in    std_logic;
    P4EL    : in    std_logic;
    P4ER    : in    std_logic;
    P4EO    : out   std_logic;
    P4RI    : in    std_logic;
    P4RL    : in    std_logic;
    P4RR    : in    std_logic;
    P4RO1   : out   std_logic;
    P4RO2   : out   std_logic;
    P4RO3   : out   std_logic;
    P4RO4   : out   std_logic;
    P4RO5   : out   std_logic;

    P5CI1   : in    std_logic;
    P5CI2   : in    std_logic;	-- DQS
    P5CI3   : in    std_logic;	-- DQS
    P5CI4   : in    std_logic;	-- DQS
    P5CI5   : in    std_logic;	-- DQS
    P5CL    : in    std_logic;
    P5CR    : in    std_logic;
    P5CO    : out   std_logic;
    P5CTI   : in    std_logic;
    P5CTO   : out   std_logic;
    P5EI1   : in    std_logic;
    P5EI2   : in    std_logic;
    P5EI3   : in    std_logic;
    P5EI4   : in    std_logic;
    P5EI5   : in    std_logic;
    P5EL    : in    std_logic;
    P5ER    : in    std_logic;
    P5EO    : out   std_logic;
    P5RI    : in    std_logic;
    P5RL    : in    std_logic;
    P5RR    : in    std_logic;
    P5RO1   : out   std_logic;
    P5RO2   : out   std_logic;
    P5RO3   : out   std_logic;
    P5RO4   : out   std_logic;
    P5RO5   : out   std_logic;

    P6CI1   : in    std_logic;
    P6CL    : in    std_logic;
    P6CR    : in    std_logic;
    P6CO    : out   std_logic;
    P6CTI   : in    std_logic;
    P6CTO   : out   std_logic;
    P6EI1   : in    std_logic;
    P6EI2   : in    std_logic;
    P6EI3   : in    std_logic;
    P6EI4   : in    std_logic;
    P6EI5   : in    std_logic;
    P6EL    : in    std_logic;
    P6ER    : in    std_logic;
    P6EO    : out   std_logic;
    P6RI    : in    std_logic;
    P6RL    : in    std_logic;
    P6RR    : in    std_logic;
    P6RO1   : out   std_logic;
    P6RO2   : out   std_logic;
    P6RO3   : out   std_logic;
    P6RO4   : out   std_logic;
    P6RO5   : out   std_logic;

    P7CI1   : in    std_logic;
    P7CL    : in    std_logic;
    P7CR    : in    std_logic;
    P7CO    : out   std_logic;
    P7CTI   : in    std_logic;
    P7CTO   : out   std_logic;
    P7EI1   : in    std_logic;
    P7EI2   : in    std_logic;
    P7EI3   : in    std_logic;
    P7EI4   : in    std_logic;
    P7EI5   : in    std_logic;
    P7EL    : in    std_logic;
    P7ER    : in    std_logic;
    P7EO    : out   std_logic;
    P7RI    : in    std_logic;
    P7RL    : in    std_logic;
    P7RR    : in    std_logic;
    P7RO1   : out   std_logic;
    P7RO2   : out   std_logic;
    P7RO3   : out   std_logic;
    P7RO4   : out   std_logic;
    P7RO5   : out   std_logic;

    P8CI1   : in    std_logic;
    P8CL    : in    std_logic;
    P8CR    : in    std_logic;
    P8CO    : out   std_logic;
    P8CTI   : in    std_logic;
    P8CTO   : out   std_logic;
    P8EI1   : in    std_logic;
    P8EI2   : in    std_logic;
    P8EI3   : in    std_logic;
    P8EI4   : in    std_logic;
    P8EI5   : in    std_logic;
    P8EL    : in    std_logic;
    P8ER    : in    std_logic;
    P8EO    : out   std_logic;
    P8RI    : in    std_logic;
    P8RL    : in    std_logic;
    P8RR    : in    std_logic;
    P8RO1   : out   std_logic;
    P8RO2   : out   std_logic;
    P8RO3   : out   std_logic;
    P8RO4   : out   std_logic;
    P8RO5   : out   std_logic;

    P9CI1   : in    std_logic;
    P9CL    : in    std_logic;
    P9CR    : in    std_logic;
    P9CO    : out   std_logic;
    P9CTI   : in    std_logic;
    P9CTO   : out   std_logic;
    P9EI1   : in    std_logic;
    P9EI2   : in    std_logic;
    P9EI3   : in    std_logic;
    P9EI4   : in    std_logic;
    P9EI5   : in    std_logic;
    P9EL    : in    std_logic;
    P9ER    : in    std_logic;
    P9EO    : out   std_logic;
    P9RI    : in    std_logic;
    P9RL    : in    std_logic;
    P9RR    : in    std_logic;
    P9RO1   : out   std_logic;
    P9RO2   : out   std_logic;
    P9RO3   : out   std_logic;
    P9RO4   : out   std_logic;
    P9RO5   : out   std_logic;

    P10CI1  : in    std_logic;
    P10CL   : in    std_logic;
    P10CR   : in    std_logic;
    P10CO   : out   std_logic;
    P10CTI  : in    std_logic;
    P10CTO  : out   std_logic;
    P10EI1  : in    std_logic;
    P10EI2  : in    std_logic;
    P10EI3  : in    std_logic;
    P10EI4  : in    std_logic;
    P10EI5  : in    std_logic;
    P10EL   : in    std_logic;
    P10ER   : in    std_logic;
    P10EO   : out   std_logic;
    P10RI   : in    std_logic;
    P10RL   : in    std_logic;
    P10RR   : in    std_logic;
    P10RO1  : out   std_logic;
    P10RO2  : out   std_logic;
    P10RO3  : out   std_logic;
    P10RO4  : out   std_logic;
    P10RO5  : out   std_logic;

    P11CI1  : in    std_logic;
    P11CL   : in    std_logic;
    P11CR   : in    std_logic;
    P11CO   : out   std_logic;
    P11CTI  : in    std_logic;
    P11CTO  : out   std_logic;
    P11EI1  : in    std_logic;
    P11EI2  : in    std_logic;
    P11EI3  : in    std_logic;
    P11EI4  : in    std_logic;
    P11EI5  : in    std_logic;
    P11EL   : in    std_logic;
    P11ER   : in    std_logic;
    P11EO   : out   std_logic;
    P11RI   : in    std_logic;
    P11RL   : in    std_logic;
    P11RR   : in    std_logic;
    P11RO1  : out   std_logic;
    P11RO2  : out   std_logic;
    P11RO3  : out   std_logic;
    P11RO4  : out   std_logic;
    P11RO5  : out   std_logic;

    P12CI1  : in    std_logic;
    P12CL   : in    std_logic;
    P12CR   : in    std_logic;
    P12CO   : out   std_logic;
    P12CTI  : in    std_logic;
    P12CTO  : out   std_logic;
    P12EI1  : in    std_logic;
    P12EI2  : in    std_logic;
    P12EI3  : in    std_logic;
    P12EI4  : in    std_logic;
    P12EI5  : in    std_logic;
    P12EL   : in    std_logic;
    P12ER   : in    std_logic;
    P12EO   : out   std_logic;
    P12RI   : in    std_logic;
    P12RL   : in    std_logic;
    P12RR   : in    std_logic;
    P12RO1  : out   std_logic;
    P12RO2  : out   std_logic;
    P12RO3  : out   std_logic;
    P12RO4  : out   std_logic;
    P12RO5  : out   std_logic;

    P13CI1  : in    std_logic;
    P13CL   : in    std_logic;
    P13CR   : in    std_logic;
    P13CO   : out   std_logic;
    P13CTI  : in    std_logic;
    P13CTO  : out   std_logic;
    P13EI1  : in    std_logic;
    P13EI2  : in    std_logic;
    P13EI3  : in    std_logic;
    P13EI4  : in    std_logic;
    P13EI5  : in    std_logic;
    P13EL   : in    std_logic;
    P13ER   : in    std_logic;
    P13EO   : out   std_logic;
    P13RI   : in    std_logic;
    P13RL   : in    std_logic;
    P13RR   : in    std_logic;
    P13RO1  : out   std_logic;
    P13RO2  : out   std_logic;
    P13RO3  : out   std_logic;
    P13RO4  : out   std_logic;
    P13RO5  : out   std_logic;

    P14CI1  : in    std_logic;
    P14CL   : in    std_logic;
    P14CR   : in    std_logic;
    P14CO   : out   std_logic;
    P14CTI  : in    std_logic;
    P14CTO  : out   std_logic;
    P14EI1  : in    std_logic;
    P14EI2  : in    std_logic;
    P14EI3  : in    std_logic;
    P14EI4  : in    std_logic;
    P14EI5  : in    std_logic;
    P14EL   : in    std_logic;
    P14ER   : in    std_logic;
    P14EO   : out   std_logic;
    P14RI   : in    std_logic;
    P14RL   : in    std_logic;
    P14RR   : in    std_logic;
    P14RO1  : out   std_logic;
    P14RO2  : out   std_logic;
    P14RO3  : out   std_logic;
    P14RO4  : out   std_logic;
    P14RO5  : out   std_logic;

    P15CI1  : in    std_logic;
    P15CL   : in    std_logic;
    P15CR   : in    std_logic;
    P15CO   : out   std_logic;
    P15CTI  : in    std_logic;
    P15CTO  : out   std_logic;
    P15EI1  : in    std_logic;
    P15EI2  : in    std_logic;
    P15EI3  : in    std_logic;
    P15EI4  : in    std_logic;
    P15EI5  : in    std_logic;
    P15EL   : in    std_logic;
    P15ER   : in    std_logic;
    P15EO   : out   std_logic;
    P15RI   : in    std_logic;
    P15RL   : in    std_logic;
    P15RR   : in    std_logic;
    P15RO1  : out   std_logic;
    P15RO2  : out   std_logic;
    P15RO3  : out   std_logic;
    P15RO4  : out   std_logic;
    P15RO5  : out   std_logic;

    P16CI1  : in    std_logic;
    P16CL   : in    std_logic;
    P16CR   : in    std_logic;
    P16CO   : out   std_logic;
    P16CTI  : in    std_logic;
    P16CTO  : out   std_logic;
    P16EI1  : in    std_logic;
    P16EI2  : in    std_logic;
    P16EI3  : in    std_logic;
    P16EI4  : in    std_logic;
    P16EI5  : in    std_logic;
    P16EL   : in    std_logic;
    P16ER   : in    std_logic;
    P16EO   : out   std_logic;
    P16RI   : in    std_logic;
    P16RL   : in    std_logic;
    P16RR   : in    std_logic;
    P16RO1  : out   std_logic;
    P16RO2  : out   std_logic;
    P16RO3  : out   std_logic;
    P16RO4  : out   std_logic;
    P16RO5  : out   std_logic;

    P17CI1  : in    std_logic;
    P17CL   : in    std_logic;
    P17CR   : in    std_logic;
    P17CO   : out   std_logic;
    P17CTI  : in    std_logic;
    P17CTO  : out   std_logic;
    P17EI1  : in    std_logic;
    P17EI2  : in    std_logic;
    P17EI3  : in    std_logic;
    P17EI4  : in    std_logic;
    P17EI5  : in    std_logic;
    P17EL   : in    std_logic;
    P17ER   : in    std_logic;
    P17EO   : out   std_logic;
    P17RI   : in    std_logic;
    P17RL   : in    std_logic;
    P17RR   : in    std_logic;
    P17RO1  : out   std_logic;
    P17RO2  : out   std_logic;
    P17RO3  : out   std_logic;
    P17RO4  : out   std_logic;
    P17RO5  : out   std_logic;

    P18CI1  : in    std_logic;
    P18CL   : in    std_logic;
    P18CR   : in    std_logic;
    P18CO   : out   std_logic;
    P18CTI  : in    std_logic;
    P18CTO  : out   std_logic;
    P18EI1  : in    std_logic;
    P18EI2  : in    std_logic;
    P18EI3  : in    std_logic;
    P18EI4  : in    std_logic;
    P18EI5  : in    std_logic;
    P18EL   : in    std_logic;
    P18ER   : in    std_logic;
    P18EO   : out   std_logic;
    P18RI   : in    std_logic;
    P18RL   : in    std_logic;
    P18RR   : in    std_logic;
    P18RO1  : out   std_logic;
    P18RO2  : out   std_logic;
    P18RO3  : out   std_logic;
    P18RO4  : out   std_logic;
    P18RO5  : out   std_logic;

    P19CI1  : in    std_logic;
    P19CL   : in    std_logic;
    P19CR   : in    std_logic;
    P19CO   : out   std_logic;
    P19CTI  : in    std_logic;
    P19CTO  : out   std_logic;
    P19EI1  : in    std_logic;
    P19EI2  : in    std_logic;
    P19EI3  : in    std_logic;
    P19EI4  : in    std_logic;
    P19EI5  : in    std_logic;
    P19EL   : in    std_logic;
    P19ER   : in    std_logic;
    P19EO   : out   std_logic;
    P19RI   : in    std_logic;
    P19RL   : in    std_logic;
    P19RR   : in    std_logic;
    P19RO1  : out   std_logic;
    P19RO2  : out   std_logic;
    P19RO3  : out   std_logic;
    P19RO4  : out   std_logic;
    P19RO5  : out   std_logic;

    P20CI1  : in    std_logic;
    P20CL   : in    std_logic;
    P20CR   : in    std_logic;
    P20CO   : out   std_logic;
    P20CTI  : in    std_logic;
    P20CTO  : out   std_logic;
    P20EI1  : in    std_logic;
    P20EI2  : in    std_logic;
    P20EI3  : in    std_logic;
    P20EI4  : in    std_logic;
    P20EI5  : in    std_logic;
    P20EL   : in    std_logic;
    P20ER   : in    std_logic;
    P20EO   : out   std_logic;
    P20RI   : in    std_logic;
    P20RL   : in    std_logic;
    P20RR   : in    std_logic;
    P20RO1  : out   std_logic;
    P20RO2  : out   std_logic;
    P20RO3  : out   std_logic;
    P20RO4  : out   std_logic;
    P20RO5  : out   std_logic;

    P21CI1  : in    std_logic;
    P21CL   : in    std_logic;
    P21CR   : in    std_logic;
    P21CO   : out   std_logic;
    P21CTI  : in    std_logic;
    P21CTO  : out   std_logic;
    P21EI1  : in    std_logic;
    P21EI2  : in    std_logic;
    P21EI3  : in    std_logic;
    P21EI4  : in    std_logic;
    P21EI5  : in    std_logic;
    P21EL   : in    std_logic;
    P21ER   : in    std_logic;
    P21EO   : out   std_logic;
    P21RI   : in    std_logic;
    P21RL   : in    std_logic;
    P21RR   : in    std_logic;
    P21RO1  : out   std_logic;
    P21RO2  : out   std_logic;
    P21RO3  : out   std_logic;
    P21RO4  : out   std_logic;
    P21RO5  : out   std_logic;

    P22CI1  : in    std_logic;
    P22CL   : in    std_logic;
    P22CR   : in    std_logic;
    P22CO   : out   std_logic;
    P22CTI  : in    std_logic;
    P22CTO  : out   std_logic;
    P22EI1  : in    std_logic;
    P22EI2  : in    std_logic;
    P22EI3  : in    std_logic;
    P22EI4  : in    std_logic;
    P22EI5  : in    std_logic;
    P22EL   : in    std_logic;
    P22ER   : in    std_logic;
    P22EO   : out   std_logic;
    P22RI   : in    std_logic;
    P22RL   : in    std_logic;
    P22RR   : in    std_logic;
    P22RO1  : out   std_logic;
    P22RO2  : out   std_logic;
    P22RO3  : out   std_logic;
    P22RO4  : out   std_logic;
    P22RO5  : out   std_logic;

    P23CI1  : in    std_logic;
    P23CL   : in    std_logic;
    P23CR   : in    std_logic;
    P23CO   : out   std_logic;
    P23CTI  : in    std_logic;
    P23CTO  : out   std_logic;
    P23EI1  : in    std_logic;
    P23EI2  : in    std_logic;
    P23EI3  : in    std_logic;
    P23EI4  : in    std_logic;
    P23EI5  : in    std_logic;
    P23EL   : in    std_logic;
    P23ER   : in    std_logic;
    P23EO   : out   std_logic;
    P23RI   : in    std_logic;
    P23RL   : in    std_logic;
    P23RR   : in    std_logic;
    P23RO1  : out   std_logic;
    P23RO2  : out   std_logic;
    P23RO3  : out   std_logic;
    P23RO4  : out   std_logic;
    P23RO5  : out   std_logic;

    P24CI1  : in    std_logic;
    P24CL   : in    std_logic;
    P24CR   : in    std_logic;
    P24CO   : out   std_logic;
    P24CTI  : in    std_logic;
    P24CTO  : out   std_logic;
    P24EI1  : in    std_logic;
    P24EI2  : in    std_logic;
    P24EI3  : in    std_logic;
    P24EI4  : in    std_logic;
    P24EI5  : in    std_logic;
    P24EL   : in    std_logic;
    P24ER   : in    std_logic;
    P24EO   : out   std_logic;
    P24RI   : in    std_logic;
    P24RL   : in    std_logic;
    P24RR   : in    std_logic;
    P24RO1  : out   std_logic;
    P24RO2  : out   std_logic;
    P24RO3  : out   std_logic;
    P24RO4  : out   std_logic;
    P24RO5  : out   std_logic;

    P25CI1  : in    std_logic;
    P25CL   : in    std_logic;
    P25CR   : in    std_logic;
    P25CO   : out   std_logic;
    P25CTI  : in    std_logic;
    P25CTO  : out   std_logic;
    P25EI1  : in    std_logic;
    P25EI2  : in    std_logic;
    P25EI3  : in    std_logic;
    P25EI4  : in    std_logic;
    P25EI5  : in    std_logic;
    P25EL   : in    std_logic;
    P25ER   : in    std_logic;
    P25EO   : out   std_logic;
    P25RI   : in    std_logic;
    P25RL   : in    std_logic;
    P25RR   : in    std_logic;
    P25RO1  : out   std_logic;
    P25RO2  : out   std_logic;
    P25RO3  : out   std_logic;
    P25RO4  : out   std_logic;
    P25RO5  : out   std_logic;

    P26CI1  : in    std_logic;
    P26CL   : in    std_logic;
    P26CR   : in    std_logic;
    P26CO   : out   std_logic;
    P26CTI  : in    std_logic;
    P26CTO  : out   std_logic;
    P26EI1  : in    std_logic;
    P26EI2  : in    std_logic;
    P26EI3  : in    std_logic;
    P26EI4  : in    std_logic;
    P26EI5  : in    std_logic;
    P26EL   : in    std_logic;
    P26ER   : in    std_logic;
    P26EO   : out   std_logic;
    P26RI   : in    std_logic;
    P26RL   : in    std_logic;
    P26RR   : in    std_logic;
    P26RO1  : out   std_logic;
    P26RO2  : out   std_logic;
    P26RO3  : out   std_logic;
    P26RO4  : out   std_logic;
    P26RO5  : out   std_logic;

    P27CI1  : in    std_logic;
    P27CL   : in    std_logic;
    P27CR   : in    std_logic;
    P27CO   : out   std_logic;
    P27CTI  : in    std_logic;
    P27CTO  : out   std_logic;
    P27EI1  : in    std_logic;
    P27EI2  : in    std_logic;
    P27EI3  : in    std_logic;
    P27EI4  : in    std_logic;
    P27EI5  : in    std_logic;
    P27EL   : in    std_logic;
    P27ER   : in    std_logic;
    P27EO   : out   std_logic;
    P27RI   : in    std_logic;
    P27RL   : in    std_logic;
    P27RR   : in    std_logic;
    P27RO1  : out   std_logic;
    P27RO2  : out   std_logic;
    P27RO3  : out   std_logic;
    P27RO4  : out   std_logic;
    P27RO5  : out   std_logic;

    P28CI1  : in    std_logic;
    P28CL   : in    std_logic;
    P28CR   : in    std_logic;
    P28CO   : out   std_logic;
    P28CTI  : in    std_logic;
    P28CTO  : out   std_logic;
    P28EI1  : in    std_logic;
    P28EI2  : in    std_logic;
    P28EI3  : in    std_logic;
    P28EI4  : in    std_logic;
    P28EI5  : in    std_logic;
    P28EL   : in    std_logic;
    P28ER   : in    std_logic;
    P28EO   : out   std_logic;
    P28RI   : in    std_logic;
    P28RL   : in    std_logic;
    P28RR   : in    std_logic;
    P28RO1  : out   std_logic;
    P28RO2  : out   std_logic;
    P28RO3  : out   std_logic;
    P28RO4  : out   std_logic;
    P28RO5  : out   std_logic;

    P29CI1  : in    std_logic;
    P29CI2  : in    std_logic;	-- DQS
    P29CI3  : in    std_logic;	-- DQS
    P29CI4  : in    std_logic;	-- DQS
    P29CI5  : in    std_logic;	-- DQS
    P29CL   : in    std_logic;
    P29CR   : in    std_logic;
    P29CO   : out   std_logic;
    P29CTI  : in    std_logic;
    P29CTO  : out   std_logic;
    P29EI1  : in    std_logic;
    P29EI2  : in    std_logic;
    P29EI3  : in    std_logic;
    P29EI4  : in    std_logic;
    P29EI5  : in    std_logic;
    P29EL   : in    std_logic;
    P29ER   : in    std_logic;
    P29EO   : out   std_logic;
    P29RI   : in    std_logic;
    P29RL   : in    std_logic;
    P29RR   : in    std_logic;
    P29RO1  : out   std_logic;
    P29RO2  : out   std_logic;
    P29RO3  : out   std_logic;
    P29RO4  : out   std_logic;
    P29RO5  : out   std_logic;

    P30CI1  : in    std_logic;
    P30CL   : in    std_logic;
    P30CR   : in    std_logic;
    P30CO   : out   std_logic;
    P30CTI  : in    std_logic;
    P30CTO  : out   std_logic;
    P30EI1  : in    std_logic;
    P30EI2  : in    std_logic;
    P30EI3  : in    std_logic;
    P30EI4  : in    std_logic;
    P30EI5  : in    std_logic;
    P30EL   : in    std_logic;
    P30ER   : in    std_logic;
    P30EO   : out   std_logic;
    P30RI   : in    std_logic;
    P30RL   : in    std_logic;
    P30RR   : in    std_logic;
    P30RO1  : out   std_logic;
    P30RO2  : out   std_logic;
    P30RO3  : out   std_logic;
    P30RO4  : out   std_logic;
    P30RO5  : out   std_logic;

    P31CI1  : in    std_logic;
    P31CL   : in    std_logic;
    P31CR   : in    std_logic;
    P31CO   : out   std_logic;
    P31CTI  : in    std_logic;
    P31CTO  : out   std_logic;
    P31EI1  : in    std_logic;
    P31EI2  : in    std_logic;
    P31EI3  : in    std_logic;
    P31EI4  : in    std_logic;
    P31EI5  : in    std_logic;
    P31EL   : in    std_logic;
    P31ER   : in    std_logic;
    P31EO   : out   std_logic;
    P31RI   : in    std_logic;
    P31RL   : in    std_logic;
    P31RR   : in    std_logic;
    P31RO1  : out   std_logic;
    P31RO2  : out   std_logic;
    P31RO3  : out   std_logic;
    P31RO4  : out   std_logic;
    P31RO5  : out   std_logic;

    P32CI1  : in    std_logic;
    P32CL   : in    std_logic;
    P32CR   : in    std_logic;
    P32CO   : out   std_logic;
    P32CTI  : in    std_logic;
    P32CTO  : out   std_logic;
    P32EI1  : in    std_logic;
    P32EI2  : in    std_logic;
    P32EI3  : in    std_logic;
    P32EI4  : in    std_logic;
    P32EI5  : in    std_logic;
    P32EL   : in    std_logic;
    P32ER   : in    std_logic;
    P32EO   : out   std_logic;
    P32RI   : in    std_logic;
    P32RL   : in    std_logic;
    P32RR   : in    std_logic;
    P32RO1  : out   std_logic;
    P32RO2  : out   std_logic;
    P32RO3  : out   std_logic;
    P32RO4  : out   std_logic;
    P32RO5  : out   std_logic;

    P33CI1  : in    std_logic;
    P33CL   : in    std_logic;
    P33CR   : in    std_logic;
    P33CO   : out   std_logic;
    P33CTI  : in    std_logic;
    P33CTO  : out   std_logic;
    P33EI1  : in    std_logic;
    P33EI2  : in    std_logic;
    P33EI3  : in    std_logic;
    P33EI4  : in    std_logic;
    P33EI5  : in    std_logic;
    P33EL   : in    std_logic;
    P33ER   : in    std_logic;
    P33EO   : out   std_logic;
    P33RI   : in    std_logic;
    P33RL   : in    std_logic;
    P33RR   : in    std_logic;
    P33RO1  : out   std_logic;
    P33RO2  : out   std_logic;
    P33RO3  : out   std_logic;
    P33RO4  : out   std_logic;
    P33RO5  : out   std_logic;

    P34CI1  : in    std_logic;
    P34CL   : in    std_logic;
    P34CR   : in    std_logic;
    P34CO   : out   std_logic;
    P34CTI  : in    std_logic;
    P34CTO  : out   std_logic;
    P34EI1  : in    std_logic;
    P34EI2  : in    std_logic;
    P34EI3  : in    std_logic;
    P34EI4  : in    std_logic;
    P34EI5  : in    std_logic;
    P34EL   : in    std_logic;
    P34ER   : in    std_logic;
    P34EO   : out   std_logic;
    P34RI   : in    std_logic;
    P34RL   : in    std_logic;
    P34RR   : in    std_logic;
    P34RO1  : out   std_logic;
    P34RO2  : out   std_logic;
    P34RO3  : out   std_logic;
    P34RO4  : out   std_logic;
    P34RO5  : out   std_logic
);
end NX_IOM_L;

-- =================================================================================================
--   NX_IOM_CONTROL_L definition                                                         2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_CONTROL_L is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port(
    RTCK1   : in    std_logic;
    RRCK1   : in    std_logic;
    WTCK1   : in    std_logic;
    WRCK1   : in    std_logic;
    RTCK2   : in    std_logic;
    RRCK2   : in    std_logic;
    WTCK2   : in    std_logic;
    WRCK2   : in    std_logic;
    CTCK    : in    std_logic;

    C1TW    : in    std_logic;
    C1TS    : in    std_logic;
    C1RW1   : in    std_logic;
    C1RW2   : in    std_logic;
    C1RW3   : in    std_logic;
    C1RNE   : in    std_logic;
    C1RS    : in    std_logic;
    C2TW    : in    std_logic;
    C2TS    : in    std_logic;
    C2RW1   : in    std_logic;
    C2RW2   : in    std_logic;
    C2RW3   : in    std_logic;
    C2RNE   : in    std_logic;
    C2RS    : in    std_logic;
    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;
    DC      : in    std_logic;
    CCK     : in    std_logic;
    DCK     : in    std_logic;
    DRI1    : in    std_logic;
    DRI2    : in    std_logic;
    DRI3    : in    std_logic;
    DRI4    : in    std_logic;
    DRI5    : in    std_logic;
    DRI6    : in    std_logic;
    DRA1    : in    std_logic;
    DRA2    : in    std_logic;
    DRA3    : in    std_logic;
    DRA4    : in    std_logic;
    DRA5    : in    std_logic;
    DRA6    : in    std_logic;
    DRL     : in    std_logic;
    DOS     : in    std_logic;
    DOG     : in    std_logic;
    DIS     : in    std_logic;
    DIG     : in    std_logic;
    DPAS    : in    std_logic;
    DPAG    : in    std_logic;
    DQSS    : in    std_logic;
    DQSG    : in    std_logic;
    DS1     : in    std_logic;
    DS2     : in    std_logic;
    CAD1    : in    std_logic;
    CAD2    : in    std_logic;
    CAD3    : in    std_logic;
    CAD4    : in    std_logic;
    CAD5    : in    std_logic;
    CAD6    : in    std_logic;
    CAP1    : in    std_logic;
    CAP2    : in    std_logic;
    CAP3    : in    std_logic;
    CAP4    : in    std_logic;
    CAN1    : in    std_logic;
    CAN2    : in    std_logic;
    CAN3    : in    std_logic;
    CAN4    : in    std_logic;
    CAT1    : in    std_logic;
    CAT2    : in    std_logic;
    CAT3    : in    std_logic;
    CAT4    : in    std_logic;
    CKO1    : out   std_logic;
    CKO2    : out   std_logic;
    FLD     : out   std_logic;
    FLG     : out   std_logic;
    C1RED   : out   std_logic;
    C2RED   : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;
    CAL     : out   std_logic;

    LINK1  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK2  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK3  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK4  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK5  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK6  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK7  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK8  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK9  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK10 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK11 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK12 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK13 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK14 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK15 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK16 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK17 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK18 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK19 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK20 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK21 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK22 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK23 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK24 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK25 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK26 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK27 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK28 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK29 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK30 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK31 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK32 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK33 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK34 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_CONTROL_L;
-- =================================================================================================
--   NX_IOM_DRIVER_M definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_DRIVER_M is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit_vector(1 downto 0) := "00";

    variant         : string := "";
    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1  : in  std_logic;
    EI2  : in  std_logic;
    EI3  : in  std_logic;
    EI4  : in  std_logic;
    EI5  : in  std_logic;
    EL   : in  std_logic;
    ER   : in  std_logic;
    CI1  : in  std_logic;
    CI2  : in  std_logic;
    CI3  : in  std_logic;
    CI4  : in  std_logic;
    CI5  : in  std_logic;
    CL   : in  std_logic;
    CR   : in  std_logic;
    CTI  : in  std_logic;
    RI   : in  std_logic;
    RL   : in  std_logic;
    RR   : in  std_logic;
    CO   : out std_logic;
    EO   : out std_logic;
    RO1  : out std_logic;
    RO2  : out std_logic;
    RO3  : out std_logic;
    RO4  : out std_logic;
    RO5  : out std_logic;
    CTO  : out std_logic;
    LINK : inout  std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_DRIVER_M;

-- =================================================================================================
--   NX_IOM_SERDES_M definition                                                          2018/10/15
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_SERDES_M is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    RTCK  : in std_logic;
    WRCK  : in std_logic;
    WTCK  : in std_logic;
    RRCK  : in std_logic;
    TRST  : in std_logic;
    RRST  : in std_logic;
    CTCK  : in std_logic;
    DCK   : in std_logic;
    DRL   : in std_logic;
    DIG   : in std_logic;
    DS    : in std_logic_vector(1 downto 0);
    DRA   : in std_logic_vector(5 downto 0);
    DRI   : in std_logic_vector(5 downto 0);
    FZ    : in std_logic;
    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0);
    FLD   : out std_logic;
    FLG   : out std_logic;
    LINKN : inout std_logic_vector(IOM_LINK_SIZE-1 downto 0);
    LINKP : inout std_logic_vector(IOM_LINK_SIZE-1 downto 0)
);
end NX_IOM_SERDES_M;
-- =================================================================================================
--   NX_IOM_DRIVER definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_DRIVER is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit_vector(1 downto 0) := "00";

    variant         : string := "";
    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1  : in  std_logic;
    EI2  : in  std_logic;
    EI3  : in  std_logic;
    EI4  : in  std_logic;
    EI5  : in  std_logic;
    EL   : in  std_logic;
    ER   : in  std_logic;
    CI1  : in  std_logic;
    CI2  : in  std_logic;
    CI3  : in  std_logic;
    CI4  : in  std_logic;
    CI5  : in  std_logic;
    CL   : in  std_logic;
    CR   : in  std_logic;
    CTI  : in  std_logic;
    RI   : in  std_logic;
    RL   : in  std_logic;
    RR   : in  std_logic;
    CO   : out std_logic;
    EO   : out std_logic;
    RO1  : out std_logic;
    RO2  : out std_logic;
    RO3  : out std_logic;
    RO4  : out std_logic;
    RO5  : out std_logic;
    CTO  : out std_logic;
    LINK : inout  std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_DRIVER;

-- =================================================================================================
--   NX_IOM_CONTROL definition                                                         2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_CONTROL is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port(
    RTCK1   : in    std_logic;
    RRCK1   : in    std_logic;
    WTCK1   : in    std_logic;
    WRCK1   : in    std_logic;
    RTCK2   : in    std_logic;
    RRCK2   : in    std_logic;
    WTCK2   : in    std_logic;
    WRCK2   : in    std_logic;
    CTCK    : in    std_logic;

    C1TW    : in    std_logic;
    C1TS    : in    std_logic;
    C1RW1   : in    std_logic;
    C1RW2   : in    std_logic;
    C1RW3   : in    std_logic;
    C1RNE   : in    std_logic;
    C1RS    : in    std_logic;
    C2TW    : in    std_logic;
    C2TS    : in    std_logic;
    C2RW1   : in    std_logic;
    C2RW2   : in    std_logic;
    C2RW3   : in    std_logic;
    C2RNE   : in    std_logic;
    C2RS    : in    std_logic;
    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;
    DC      : in    std_logic;
    CCK     : in    std_logic;
    DCK     : in    std_logic;
    DRI1    : in    std_logic;
    DRI2    : in    std_logic;
    DRI3    : in    std_logic;
    DRI4    : in    std_logic;
    DRI5    : in    std_logic;
    DRI6    : in    std_logic;
    DRA1    : in    std_logic;
    DRA2    : in    std_logic;
    DRA3    : in    std_logic;
    DRA4    : in    std_logic;
    DRA5    : in    std_logic;
    DRA6    : in    std_logic;
    DRL     : in    std_logic;
    DOS     : in    std_logic;
    DOG     : in    std_logic;
    DIS     : in    std_logic;
    DIG     : in    std_logic;
    DPAS    : in    std_logic;
    DPAG    : in    std_logic;
    DQSS    : in    std_logic;
    DQSG    : in    std_logic;
    DS1     : in    std_logic;
    DS2     : in    std_logic;
    CAD1    : in    std_logic;
    CAD2    : in    std_logic;
    CAD3    : in    std_logic;
    CAD4    : in    std_logic;
    CAD5    : in    std_logic;
    CAD6    : in    std_logic;
    CAP1    : in    std_logic;
    CAP2    : in    std_logic;
    CAP3    : in    std_logic;
    CAP4    : in    std_logic;
    CAN1    : in    std_logic;
    CAN2    : in    std_logic;
    CAN3    : in    std_logic;
    CAN4    : in    std_logic;
    CAT1    : in    std_logic;
    CAT2    : in    std_logic;
    CAT3    : in    std_logic;
    CAT4    : in    std_logic;
    SPI1    : in    std_logic;
    SPI2    : in    std_logic;
    SPI3    : in    std_logic;
    CKO1    : out   std_logic;
    CKO2    : out   std_logic;
    FLD     : out   std_logic;
    FLG     : out   std_logic;
    C1RED   : out   std_logic;
    C2RED   : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;
    CAL     : out   std_logic;

    LINK1  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK2  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK3  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK4  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK5  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK6  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK7  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK8  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK9  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK10 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK11 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK12 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK13 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK14 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK15 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK16 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK17 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK18 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK19 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK20 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK21 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK22 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK23 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK24 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK25 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK26 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK27 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK28 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK29 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK30 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK31 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK32 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK33 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK34 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_CONTROL;

-- =================================================================================================
--   NX_IOM_SERDES definition                                                          2018/10/15
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_SERDES is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    RTCK  : in std_logic;
    WRCK  : in std_logic;
    WTCK  : in std_logic;
    RRCK  : in std_logic;
    TRST  : in std_logic;
    RRST  : in std_logic;
    CTCK  : in std_logic;
    DCK   : in std_logic;
    DRL   : in std_logic;
    DIG   : in std_logic;
    DS    : in std_logic_vector(1 downto 0);
    DRA   : in std_logic_vector(5 downto 0);
    DRI   : in std_logic_vector(5 downto 0);
    FZ    : in std_logic;
    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0);
    FLD   : out std_logic;
    FLG   : out std_logic;
    LINKN : inout std_logic_vector(IOM_LINK_SIZE-1 downto 0);
    LINKP : inout std_logic_vector(IOM_LINK_SIZE-1 downto 0)
);
end NX_IOM_SERDES;

-- =================================================================================================
--   Wrappers to new name
-- =================================================================================================

--NX_IOM_DRIVER##{{{##
architecture NX_RTL of NX_IOM_DRIVER is
begin

    process (CTI) begin				-- Dummy input for syntax analysis
	report "Model NX_IOM_DRIVER is superceded by NX_IOM_DRIVER_M" severity note;
    end process;


base : NX_IOM_DRIVER_M
generic map (
    epath_edge     => epath_edge,
    epath_init     => epath_init,
    epath_load     => epath_load,
    epath_mode     => epath_mode,
    epath_sync     => epath_sync,
    epath_dynamic  => epath_dynamic,

    rpath_edge     => rpath_edge,
    rpath_init     => rpath_init,
    rpath_load     => rpath_load,
    rpath_mode     => rpath_mode,
    rpath_sync     => rpath_sync,
    rpath_dynamic  => rpath_dynamic,

    cpath_edge     => cpath_edge,
    cpath_init     => cpath_init,
    cpath_load     => cpath_load,
    cpath_mode     => cpath_mode,
    cpath_sync     => cpath_sync,
    cpath_inv      => cpath_inv,

    tpath_mode     => tpath_mode,

    variant        => variant,
    location       => location,
    chained        => chained,
    symbol         => symbol
)
port map (
    EI1  => EI1,
    EI2  => EI2,
    EI3  => EI3,
    EI4  => EI4,
    EI5  => EI5,
    EL   => EL,
    ER   => ER,
    CI1  => CI1,
    CI2  => CI2,
    CI3  => CI3,
    CI4  => CI4,
    CI5  => CI5,
    CL   => CL,
    CR   => CR,
    CTI  => CTI,
    RI   => RI,
    RL   => RL,
    RR   => RR,
    CO   => CO,
    EO   => EO,
    RO1  => RO1,
    RO2  => RO2,
    RO3  => RO3,
    RO4  => RO4,
    RO5  => RO5,
    CTO  => CTO,
    LINK => LINK
);

end NX_RTL;
--##}}}##

--NX_IOM_CONTROL##{{{##
architecture NX_RTL of NX_IOM_CONTROL is
begin

    process (CTCK) begin			-- Dummy input for syntax analysis
	report "Model NX_IOM_CONTROL is superceded by NX_IOM_CONTROL_M" severity note;
    end process;

base : NX_IOM_CONTROL_M
generic map (
    mode_side1   => mode_side1,
    sel_clkw_rx1 => sel_clkw_rx1,
    sel_clkr_rx1 => sel_clkr_rx1,
    div_tx1      => div_tx1,
    div_rx1      => div_rx1,
    inv_di_fclk1 => inv_di_fclk1,
    latency1     => latency1,
    mode_side2   => mode_side2,
    sel_clkw_rx2 => sel_clkw_rx2,
    sel_clkr_rx2 => sel_clkr_rx2,
    div_tx2      => div_tx2,
    div_rx2      => div_rx2,
    inv_di_fclk2 => inv_di_fclk2,
    latency2     => latency2,
    sel_clk_out1 => sel_clk_out1,
    sel_clk_out2 => sel_clk_out2,
    mode_rpath   => mode_rpath,
    mode_epath   => mode_epath,
    mode_cpath   => mode_cpath,
    mode_tpath   => mode_tpath,
    mode_io_cal  => mode_io_cal,
    location     => location
)
port map (
    RTCK1  => RTCK1,
    RRCK1  => RRCK1,
    WTCK1  => WTCK1,
    WRCK1  => WRCK1,
    RTCK2  => RTCK2,
    RRCK2  => RRCK2,
    WTCK2  => WTCK2,
    WRCK2  => WRCK2,
    CTCK   => CTCK,

    C1TW   => C1TW,
    C1TS   => C1TS,
    C1RW1  => C1RW1,
    C1RW2  => C1RW2,
    C1RW3  => C1RW3,
    C1RNE  => C1RNE,
    C1RS   => C1RS,
    C2TW   => C2TW,
    C2TS   => C2TS,
    C2RW1  => C2RW1,
    C2RW2  => C2RW2,
    C2RW3  => C2RW3,
    C2RNE  => C2RNE,
    C2RS   => C2RS,
    FA1    => FA1,
    FA2    => FA2,
    FA3    => FA3,
    FA4    => FA4,
    FA5    => FA5,
    FA6    => FA6,
    FZ     => FZ,
    DC     => DC,
    CCK    => CCK,
    DCK    => DCK,
    DRI1   => DRI1,
    DRI2   => DRI2,
    DRI3   => DRI3,
    DRI4   => DRI4,
    DRI5   => DRI5,
    DRI6   => DRI6,
    DRA1   => DRA1,
    DRA2   => DRA2,
    DRA3   => DRA3,
    DRA4   => DRA4,
    DRA5   => DRA5,
    DRA6   => DRA6,
    DRL    => DRL,
    DOS    => DOS,
    DOG    => DOG,
    DIS    => DIS,
    DIG    => DIG,
    DPAS   => DPAS,
    DPAG   => DPAG,
    DQSS   => DQSS,
    DQSG   => DQSG,
    DS1    => DS1,
    DS2    => DS2,
    CAD1   => CAD1,
    CAD2   => CAD2,
    CAD3   => CAD3,
    CAD4   => CAD4,
    CAD5   => CAD5,
    CAD6   => CAD6,
    CAP1   => CAP1,
    CAP2   => CAP2,
    CAP3   => CAP3,
    CAP4   => CAP4,
    CAN1   => CAN1,
    CAN2   => CAN2,
    CAN3   => CAN3,
    CAN4   => CAN4,
    CAT1   => CAT1,
    CAT2   => CAT2,
    CAT3   => CAT3,
    CAT4   => CAT4,
    SPI1   => SPI1,
    SPI2   => SPI2,
    SPI3   => SPI3,
    CKO1   => CKO1,
    CKO2   => CKO2,
    FLD    => FLD,
    FLG    => FLG,
    C1RED  => C1RED,
    C2RED  => C2RED,
    DRO1   => DRO1,
    DRO2   => DRO2,
    DRO3   => DRO3,
    DRO4   => DRO4,
    DRO5   => DRO5,
    DRO6   => DRO6,
    CAL    => CAL,

    LINK1  => LINK1,
    LINK2  => LINK2,
    LINK3  => LINK3,
    LINK4  => LINK4,
    LINK5  => LINK5,
    LINK6  => LINK6,
    LINK7  => LINK7,
    LINK8  => LINK8,
    LINK9  => LINK9,
    LINK10 => LINK10,
    LINK11 => LINK11,
    LINK12 => LINK12,
    LINK13 => LINK13,
    LINK14 => LINK14,
    LINK15 => LINK15,
    LINK16 => LINK16,
    LINK17 => LINK17,
    LINK18 => LINK18,
    LINK19 => LINK19,
    LINK20 => LINK20,
    LINK21 => LINK21,
    LINK22 => LINK22,
    LINK23 => LINK23,
    LINK24 => LINK24,
    LINK25 => LINK25,
    LINK26 => LINK26,
    LINK27 => LINK27,
    LINK28 => LINK28,
    LINK29 => LINK29,
    LINK30 => LINK30,
    LINK31 => LINK31,
    LINK32 => LINK32,
    LINK33 => LINK33,
    LINK34 => LINK34
);

end NX_RTL;
--##}}}##

--NX_IOM_SERDES##{{{##
architecture NX_RTL of NX_IOM_SERDES is
begin

    process (RTCK) begin			-- Dummy input for syntax analysis
	report "Model NX_IOM_SERDES is superceded by NX_IOM_SERDES_M" severity note;
    end process;

base : NX_IOM_SERDES_M
generic map (
    data_size => data_size,
    location  => location 
)
port map (
    RTCK  => RTCK,
    WRCK  => WRCK,
    WTCK  => WTCK,
    RRCK  => RRCK,
    TRST  => TRST,
    RRST  => RRST,
    CTCK  => CTCK,
    DCK   => DCK,
    DRL   => DRL,
    DIG   => DIG,
    DS    => DS,
    DRA   => DRA,
    DRI   => DRI,
    FZ    => FZ,
    DRO   => DRO,
    DID   => DID,
    FLD   => FLD,
    FLG   => FLG,
    LINKN => LINKN,
    LINKP => LINKP
);

end NX_RTL;
--##}}}##
-- =================================================================================================
--   NX_IOM definition                                                                  2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk1 : bit := '0';
--  latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
--  inv_di_fclk2 : bit := '0';
--  latency2     : bit := '0';
--  sel_clk_out2 : bit_vector(1 downto 0) := "00";
--  sel_clk_out3 : bit_vector(1 downto 0) := "00";
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_io_cal  : bit := '0';
    pads_dict    : string := "";
    pads_path    : string := ""
);
port(
    RTCK1   : in    std_logic;
    RRCK1   : in    std_logic;
    WTCK1   : in    std_logic;
    WRCK1   : in    std_logic;
    RTCK2   : in    std_logic;
    RRCK2   : in    std_logic;
    WTCK2   : in    std_logic;
    WRCK2   : in    std_logic;
    CTCK    : in    std_logic;
    CCK     : in    std_logic;
    DCK     : in    std_logic;

    C1TW    : in    std_logic;
    C1TS    : in    std_logic;
    C1RW1   : in    std_logic;
    C1RW2   : in    std_logic;
    C1RW3   : in    std_logic;
    C1RNE   : in    std_logic;
    C1RS    : in    std_logic;
    C2TW    : in    std_logic;
    C2TS    : in    std_logic;
    C2RW1   : in    std_logic;
    C2RW2   : in    std_logic;
    C2RW3   : in    std_logic;
    C2RNE   : in    std_logic;
    C2RS    : in    std_logic;
    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FZ      : in    std_logic;
    DC      : in    std_logic;
    DRI1    : in    std_logic;
    DRI2    : in    std_logic;
    DRI3    : in    std_logic;
    DRI4    : in    std_logic;
    DRI5    : in    std_logic;
    DRI6    : in    std_logic;
    DRA1    : in    std_logic;
    DRA2    : in    std_logic;
    DRA3    : in    std_logic;
    DRA4    : in    std_logic;
    DRA5    : in    std_logic;
    DRL     : in    std_logic;
    DOS     : in    std_logic;
    DOG     : in    std_logic;
    DIS     : in    std_logic;
    DIG     : in    std_logic;
    DPAS    : in    std_logic;
    DPAG    : in    std_logic;
    DQSS    : in    std_logic;
    DQSG    : in    std_logic;
    DS1     : in    std_logic;
    DS2     : in    std_logic;
    CAD1    : in    std_logic;
    CAD2    : in    std_logic;
    CAD3    : in    std_logic;
    CAD4    : in    std_logic;
    CAD5    : in    std_logic;
    CAD6    : in    std_logic;
    CAP1    : in    std_logic;
    CAP2    : in    std_logic;
    CAP3    : in    std_logic;
    CAP4    : in    std_logic;
    CAN1    : in    std_logic;
    CAN2    : in    std_logic;
    CAN3    : in    std_logic;
    CAN4    : in    std_logic;
    CAT1    : in    std_logic;
    CAT2    : in    std_logic;
    CAT3    : in    std_logic;
    CAT4    : in    std_logic;
    SPI1    : in    std_logic;
    SPI2    : in    std_logic;
    SPI3    : in    std_logic;

    CKO1    : out   std_logic;
    CKO2    : out   std_logic;

    FLD     : out   std_logic;
    FLG     : out   std_logic;
    C1RED   : out   std_logic;
    C2RED   : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;
    CAL     : out   std_logic;

    P1CI1   : in    std_logic;
    P1CL    : in    std_logic;
    P1CR    : in    std_logic;
    P1CO    : out   std_logic;
    P1CTI   : in    std_logic;
    P1CTO   : out   std_logic;
    P1EI1   : in    std_logic;
    P1EI2   : in    std_logic;
    P1EI3   : in    std_logic;
    P1EI4   : in    std_logic;
    P1EI5   : in    std_logic;
    P1EL    : in    std_logic;
    P1ER    : in    std_logic;
    P1EO    : out   std_logic;
    P1RI    : in    std_logic;
    P1RL    : in    std_logic;
    P1RR    : in    std_logic;
    P1RO1   : out   std_logic;
    P1RO2   : out   std_logic;
    P1RO3   : out   std_logic;
    P1RO4   : out   std_logic;
    P1RO5   : out   std_logic;

    P2CI1   : in    std_logic;
    P2CL    : in    std_logic;
    P2CR    : in    std_logic;
    P2CO    : out   std_logic;
    P2CTI   : in    std_logic;
    P2CTO   : out   std_logic;
    P2EI1   : in    std_logic;
    P2EI2   : in    std_logic;
    P2EI3   : in    std_logic;
    P2EI4   : in    std_logic;
    P2EI5   : in    std_logic;
    P2EL    : in    std_logic;
    P2ER    : in    std_logic;
    P2EO    : out   std_logic;
    P2RI    : in    std_logic;
    P2RL    : in    std_logic;
    P2RR    : in    std_logic;
    P2RO1   : out   std_logic;
    P2RO2   : out   std_logic;
    P2RO3   : out   std_logic;
    P2RO4   : out   std_logic;
    P2RO5   : out   std_logic;

    P3CI1   : in    std_logic;
    P3CL    : in    std_logic;
    P3CR    : in    std_logic;
    P3CO    : out   std_logic;
    P3CTI   : in    std_logic;
    P3CTO   : out   std_logic;
    P3EI1   : in    std_logic;
    P3EI2   : in    std_logic;
    P3EI3   : in    std_logic;
    P3EI4   : in    std_logic;
    P3EI5   : in    std_logic;
    P3EL    : in    std_logic;
    P3ER    : in    std_logic;
    P3EO    : out   std_logic;
    P3RI    : in    std_logic;
    P3RL    : in    std_logic;
    P3RR    : in    std_logic;
    P3RO1   : out   std_logic;
    P3RO2   : out   std_logic;
    P3RO3   : out   std_logic;
    P3RO4   : out   std_logic;
    P3RO5   : out   std_logic;

    P4CI1   : in    std_logic;
    P4CL    : in    std_logic;
    P4CR    : in    std_logic;
    P4CO    : out   std_logic;
    P4CTI   : in    std_logic;
    P4CTO   : out   std_logic;
    P4EI1   : in    std_logic;
    P4EI2   : in    std_logic;
    P4EI3   : in    std_logic;
    P4EI4   : in    std_logic;
    P4EI5   : in    std_logic;
    P4EL    : in    std_logic;
    P4ER    : in    std_logic;
    P4EO    : out   std_logic;
    P4RI    : in    std_logic;
    P4RL    : in    std_logic;
    P4RR    : in    std_logic;
    P4RO1   : out   std_logic;
    P4RO2   : out   std_logic;
    P4RO3   : out   std_logic;
    P4RO4   : out   std_logic;
    P4RO5   : out   std_logic;

    P5CI1   : in    std_logic;
    P5CI2   : in    std_logic;	-- DQS
    P5CI3   : in    std_logic;	-- DQS
    P5CI4   : in    std_logic;	-- DQS
    P5CI5   : in    std_logic;	-- DQS
    P5CL    : in    std_logic;
    P5CR    : in    std_logic;
    P5CO    : out   std_logic;
    P5CTI   : in    std_logic;
    P5CTO   : out   std_logic;
    P5EI1   : in    std_logic;
    P5EI2   : in    std_logic;
    P5EI3   : in    std_logic;
    P5EI4   : in    std_logic;
    P5EI5   : in    std_logic;
    P5EL    : in    std_logic;
    P5ER    : in    std_logic;
    P5EO    : out   std_logic;
    P5RI    : in    std_logic;
    P5RL    : in    std_logic;
    P5RR    : in    std_logic;
    P5RO1   : out   std_logic;
    P5RO2   : out   std_logic;
    P5RO3   : out   std_logic;
    P5RO4   : out   std_logic;
    P5RO5   : out   std_logic;

    P6CI1   : in    std_logic;
    P6CL    : in    std_logic;
    P6CR    : in    std_logic;
    P6CO    : out   std_logic;
    P6CTI   : in    std_logic;
    P6CTO   : out   std_logic;
    P6EI1   : in    std_logic;
    P6EI2   : in    std_logic;
    P6EI3   : in    std_logic;
    P6EI4   : in    std_logic;
    P6EI5   : in    std_logic;
    P6EL    : in    std_logic;
    P6ER    : in    std_logic;
    P6EO    : out   std_logic;
    P6RI    : in    std_logic;
    P6RL    : in    std_logic;
    P6RR    : in    std_logic;
    P6RO1   : out   std_logic;
    P6RO2   : out   std_logic;
    P6RO3   : out   std_logic;
    P6RO4   : out   std_logic;
    P6RO5   : out   std_logic;

    P7CI1   : in    std_logic;
    P7CL    : in    std_logic;
    P7CR    : in    std_logic;
    P7CO    : out   std_logic;
    P7CTI   : in    std_logic;
    P7CTO   : out   std_logic;
    P7EI1   : in    std_logic;
    P7EI2   : in    std_logic;
    P7EI3   : in    std_logic;
    P7EI4   : in    std_logic;
    P7EI5   : in    std_logic;
    P7EL    : in    std_logic;
    P7ER    : in    std_logic;
    P7EO    : out   std_logic;
    P7RI    : in    std_logic;
    P7RL    : in    std_logic;
    P7RR    : in    std_logic;
    P7RO1   : out   std_logic;
    P7RO2   : out   std_logic;
    P7RO3   : out   std_logic;
    P7RO4   : out   std_logic;
    P7RO5   : out   std_logic;

    P8CI1   : in    std_logic;
    P8CL    : in    std_logic;
    P8CR    : in    std_logic;
    P8CO    : out   std_logic;
    P8CTI   : in    std_logic;
    P8CTO   : out   std_logic;
    P8EI1   : in    std_logic;
    P8EI2   : in    std_logic;
    P8EI3   : in    std_logic;
    P8EI4   : in    std_logic;
    P8EI5   : in    std_logic;
    P8EL    : in    std_logic;
    P8ER    : in    std_logic;
    P8EO    : out   std_logic;
    P8RI    : in    std_logic;
    P8RL    : in    std_logic;
    P8RR    : in    std_logic;
    P8RO1   : out   std_logic;
    P8RO2   : out   std_logic;
    P8RO3   : out   std_logic;
    P8RO4   : out   std_logic;
    P8RO5   : out   std_logic;

    P9CI1   : in    std_logic;
    P9CL    : in    std_logic;
    P9CR    : in    std_logic;
    P9CO    : out   std_logic;
    P9CTI   : in    std_logic;
    P9CTO   : out   std_logic;
    P9EI1   : in    std_logic;
    P9EI2   : in    std_logic;
    P9EI3   : in    std_logic;
    P9EI4   : in    std_logic;
    P9EI5   : in    std_logic;
    P9EL    : in    std_logic;
    P9ER    : in    std_logic;
    P9EO    : out   std_logic;
    P9RI    : in    std_logic;
    P9RL    : in    std_logic;
    P9RR    : in    std_logic;
    P9RO1   : out   std_logic;
    P9RO2   : out   std_logic;
    P9RO3   : out   std_logic;
    P9RO4   : out   std_logic;
    P9RO5   : out   std_logic;

    P10CI1  : in    std_logic;
    P10CL   : in    std_logic;
    P10CR   : in    std_logic;
    P10CO   : out   std_logic;
    P10CTI  : in    std_logic;
    P10CTO  : out   std_logic;
    P10EI1  : in    std_logic;
    P10EI2  : in    std_logic;
    P10EI3  : in    std_logic;
    P10EI4  : in    std_logic;
    P10EI5  : in    std_logic;
    P10EL   : in    std_logic;
    P10ER   : in    std_logic;
    P10EO   : out   std_logic;
    P10RI   : in    std_logic;
    P10RL   : in    std_logic;
    P10RR   : in    std_logic;
    P10RO1  : out   std_logic;
    P10RO2  : out   std_logic;
    P10RO3  : out   std_logic;
    P10RO4  : out   std_logic;
    P10RO5  : out   std_logic;

    P11CI1  : in    std_logic;
    P11CL   : in    std_logic;
    P11CR   : in    std_logic;
    P11CO   : out   std_logic;
    P11CTI  : in    std_logic;
    P11CTO  : out   std_logic;
    P11EI1  : in    std_logic;
    P11EI2  : in    std_logic;
    P11EI3  : in    std_logic;
    P11EI4  : in    std_logic;
    P11EI5  : in    std_logic;
    P11EL   : in    std_logic;
    P11ER   : in    std_logic;
    P11EO   : out   std_logic;
    P11RI   : in    std_logic;
    P11RL   : in    std_logic;
    P11RR   : in    std_logic;
    P11RO1  : out   std_logic;
    P11RO2  : out   std_logic;
    P11RO3  : out   std_logic;
    P11RO4  : out   std_logic;
    P11RO5  : out   std_logic;

    P12CI1  : in    std_logic;
    P12CL   : in    std_logic;
    P12CR   : in    std_logic;
    P12CO   : out   std_logic;
    P12CTI  : in    std_logic;
    P12CTO  : out   std_logic;
    P12EI1  : in    std_logic;
    P12EI2  : in    std_logic;
    P12EI3  : in    std_logic;
    P12EI4  : in    std_logic;
    P12EI5  : in    std_logic;
    P12EL   : in    std_logic;
    P12ER   : in    std_logic;
    P12EO   : out   std_logic;
    P12RI   : in    std_logic;
    P12RL   : in    std_logic;
    P12RR   : in    std_logic;
    P12RO1  : out   std_logic;
    P12RO2  : out   std_logic;
    P12RO3  : out   std_logic;
    P12RO4  : out   std_logic;
    P12RO5  : out   std_logic;

    P13CI1  : in    std_logic;
    P13CL   : in    std_logic;
    P13CR   : in    std_logic;
    P13CO   : out   std_logic;
    P13CTI  : in    std_logic;
    P13CTO  : out   std_logic;
    P13EI1  : in    std_logic;
    P13EI2  : in    std_logic;
    P13EI3  : in    std_logic;
    P13EI4  : in    std_logic;
    P13EI5  : in    std_logic;
    P13EL   : in    std_logic;
    P13ER   : in    std_logic;
    P13EO   : out   std_logic;
    P13RI   : in    std_logic;
    P13RL   : in    std_logic;
    P13RR   : in    std_logic;
    P13RO1  : out   std_logic;
    P13RO2  : out   std_logic;
    P13RO3  : out   std_logic;
    P13RO4  : out   std_logic;
    P13RO5  : out   std_logic;

    P14CI1  : in    std_logic;
    P14CL   : in    std_logic;
    P14CR   : in    std_logic;
    P14CO   : out   std_logic;
    P14CTI  : in    std_logic;
    P14CTO  : out   std_logic;
    P14EI1  : in    std_logic;
    P14EI2  : in    std_logic;
    P14EI3  : in    std_logic;
    P14EI4  : in    std_logic;
    P14EI5  : in    std_logic;
    P14EL   : in    std_logic;
    P14ER   : in    std_logic;
    P14EO   : out   std_logic;
    P14RI   : in    std_logic;
    P14RL   : in    std_logic;
    P14RR   : in    std_logic;
    P14RO1  : out   std_logic;
    P14RO2  : out   std_logic;
    P14RO3  : out   std_logic;
    P14RO4  : out   std_logic;
    P14RO5  : out   std_logic;

    P15CI1  : in    std_logic;
    P15CL   : in    std_logic;
    P15CR   : in    std_logic;
    P15CO   : out   std_logic;
    P15CTI  : in    std_logic;
    P15CTO  : out   std_logic;
    P15EI1  : in    std_logic;
    P15EI2  : in    std_logic;
    P15EI3  : in    std_logic;
    P15EI4  : in    std_logic;
    P15EI5  : in    std_logic;
    P15EL   : in    std_logic;
    P15ER   : in    std_logic;
    P15EO   : out   std_logic;
    P15RI   : in    std_logic;
    P15RL   : in    std_logic;
    P15RR   : in    std_logic;
    P15RO1  : out   std_logic;
    P15RO2  : out   std_logic;
    P15RO3  : out   std_logic;
    P15RO4  : out   std_logic;
    P15RO5  : out   std_logic;

    P16CI1  : in    std_logic;
    P16CL   : in    std_logic;
    P16CR   : in    std_logic;
    P16CO   : out   std_logic;
    P16CTI  : in    std_logic;
    P16CTO  : out   std_logic;
    P16EI1  : in    std_logic;
    P16EI2  : in    std_logic;
    P16EI3  : in    std_logic;
    P16EI4  : in    std_logic;
    P16EI5  : in    std_logic;
    P16EL   : in    std_logic;
    P16ER   : in    std_logic;
    P16EO   : out   std_logic;
    P16RI   : in    std_logic;
    P16RL   : in    std_logic;
    P16RR   : in    std_logic;
    P16RO1  : out   std_logic;
    P16RO2  : out   std_logic;
    P16RO3  : out   std_logic;
    P16RO4  : out   std_logic;
    P16RO5  : out   std_logic;

    P17CI1  : in    std_logic;
    P17CL   : in    std_logic;
    P17CR   : in    std_logic;
    P17CO   : out   std_logic;
    P17CTI  : in    std_logic;
    P17CTO  : out   std_logic;
    P17EI1  : in    std_logic;
    P17EI2  : in    std_logic;
    P17EI3  : in    std_logic;
    P17EI4  : in    std_logic;
    P17EI5  : in    std_logic;
    P17EL   : in    std_logic;
    P17ER   : in    std_logic;
    P17EO   : out   std_logic;
    P17RI   : in    std_logic;
    P17RL   : in    std_logic;
    P17RR   : in    std_logic;
    P17RO1  : out   std_logic;
    P17RO2  : out   std_logic;
    P17RO3  : out   std_logic;
    P17RO4  : out   std_logic;
    P17RO5  : out   std_logic;

    P18CI1  : in    std_logic;
    P18CL   : in    std_logic;
    P18CR   : in    std_logic;
    P18CO   : out   std_logic;
    P18CTI  : in    std_logic;
    P18CTO  : out   std_logic;
    P18EI1  : in    std_logic;
    P18EI2  : in    std_logic;
    P18EI3  : in    std_logic;
    P18EI4  : in    std_logic;
    P18EI5  : in    std_logic;
    P18EL   : in    std_logic;
    P18ER   : in    std_logic;
    P18EO   : out   std_logic;
    P18RI   : in    std_logic;
    P18RL   : in    std_logic;
    P18RR   : in    std_logic;
    P18RO1  : out   std_logic;
    P18RO2  : out   std_logic;
    P18RO3  : out   std_logic;
    P18RO4  : out   std_logic;
    P18RO5  : out   std_logic;

    P19CI1  : in    std_logic;
    P19CL   : in    std_logic;
    P19CR   : in    std_logic;
    P19CO   : out   std_logic;
    P19CTI  : in    std_logic;
    P19CTO  : out   std_logic;
    P19EI1  : in    std_logic;
    P19EI2  : in    std_logic;
    P19EI3  : in    std_logic;
    P19EI4  : in    std_logic;
    P19EI5  : in    std_logic;
    P19EL   : in    std_logic;
    P19ER   : in    std_logic;
    P19EO   : out   std_logic;
    P19RI   : in    std_logic;
    P19RL   : in    std_logic;
    P19RR   : in    std_logic;
    P19RO1  : out   std_logic;
    P19RO2  : out   std_logic;
    P19RO3  : out   std_logic;
    P19RO4  : out   std_logic;
    P19RO5  : out   std_logic;

    P20CI1  : in    std_logic;
    P20CL   : in    std_logic;
    P20CR   : in    std_logic;
    P20CO   : out   std_logic;
    P20CTI  : in    std_logic;
    P20CTO  : out   std_logic;
    P20EI1  : in    std_logic;
    P20EI2  : in    std_logic;
    P20EI3  : in    std_logic;
    P20EI4  : in    std_logic;
    P20EI5  : in    std_logic;
    P20EL   : in    std_logic;
    P20ER   : in    std_logic;
    P20EO   : out   std_logic;
    P20RI   : in    std_logic;
    P20RL   : in    std_logic;
    P20RR   : in    std_logic;
    P20RO1  : out   std_logic;
    P20RO2  : out   std_logic;
    P20RO3  : out   std_logic;
    P20RO4  : out   std_logic;
    P20RO5  : out   std_logic;

    P21CI1  : in    std_logic;
    P21CL   : in    std_logic;
    P21CR   : in    std_logic;
    P21CO   : out   std_logic;
    P21CTI  : in    std_logic;
    P21CTO  : out   std_logic;
    P21EI1  : in    std_logic;
    P21EI2  : in    std_logic;
    P21EI3  : in    std_logic;
    P21EI4  : in    std_logic;
    P21EI5  : in    std_logic;
    P21EL   : in    std_logic;
    P21ER   : in    std_logic;
    P21EO   : out   std_logic;
    P21RI   : in    std_logic;
    P21RL   : in    std_logic;
    P21RR   : in    std_logic;
    P21RO1  : out   std_logic;
    P21RO2  : out   std_logic;
    P21RO3  : out   std_logic;
    P21RO4  : out   std_logic;
    P21RO5  : out   std_logic;

    P22CI1  : in    std_logic;
    P22CL   : in    std_logic;
    P22CR   : in    std_logic;
    P22CO   : out   std_logic;
    P22CTI  : in    std_logic;
    P22CTO  : out   std_logic;
    P22EI1  : in    std_logic;
    P22EI2  : in    std_logic;
    P22EI3  : in    std_logic;
    P22EI4  : in    std_logic;
    P22EI5  : in    std_logic;
    P22EL   : in    std_logic;
    P22ER   : in    std_logic;
    P22EO   : out   std_logic;
    P22RI   : in    std_logic;
    P22RL   : in    std_logic;
    P22RR   : in    std_logic;
    P22RO1  : out   std_logic;
    P22RO2  : out   std_logic;
    P22RO3  : out   std_logic;
    P22RO4  : out   std_logic;
    P22RO5  : out   std_logic;

    P23CI1  : in    std_logic;
    P23CL   : in    std_logic;
    P23CR   : in    std_logic;
    P23CO   : out   std_logic;
    P23CTI  : in    std_logic;
    P23CTO  : out   std_logic;
    P23EI1  : in    std_logic;
    P23EI2  : in    std_logic;
    P23EI3  : in    std_logic;
    P23EI4  : in    std_logic;
    P23EI5  : in    std_logic;
    P23EL   : in    std_logic;
    P23ER   : in    std_logic;
    P23EO   : out   std_logic;
    P23RI   : in    std_logic;
    P23RL   : in    std_logic;
    P23RR   : in    std_logic;
    P23RO1  : out   std_logic;
    P23RO2  : out   std_logic;
    P23RO3  : out   std_logic;
    P23RO4  : out   std_logic;
    P23RO5  : out   std_logic;

    P24CI1  : in    std_logic;
    P24CL   : in    std_logic;
    P24CR   : in    std_logic;
    P24CO   : out   std_logic;
    P24CTI  : in    std_logic;
    P24CTO  : out   std_logic;
    P24EI1  : in    std_logic;
    P24EI2  : in    std_logic;
    P24EI3  : in    std_logic;
    P24EI4  : in    std_logic;
    P24EI5  : in    std_logic;
    P24EL   : in    std_logic;
    P24ER   : in    std_logic;
    P24EO   : out   std_logic;
    P24RI   : in    std_logic;
    P24RL   : in    std_logic;
    P24RR   : in    std_logic;
    P24RO1  : out   std_logic;
    P24RO2  : out   std_logic;
    P24RO3  : out   std_logic;
    P24RO4  : out   std_logic;
    P24RO5  : out   std_logic;

    P25CI1  : in    std_logic;
    P25CI2  : in    std_logic;	-- DQS
    P25CI3  : in    std_logic;	-- DQS
    P25CI4  : in    std_logic;	-- DQS
    P25CI5  : in    std_logic;	-- DQS
    P25CL   : in    std_logic;
    P25CR   : in    std_logic;
    P25CO   : out   std_logic;
    P25CTI  : in    std_logic;
    P25CTO  : out   std_logic;
    P25EI1  : in    std_logic;
    P25EI2  : in    std_logic;
    P25EI3  : in    std_logic;
    P25EI4  : in    std_logic;
    P25EI5  : in    std_logic;
    P25EL   : in    std_logic;
    P25ER   : in    std_logic;
    P25EO   : out   std_logic;
    P25RI   : in    std_logic;
    P25RL   : in    std_logic;
    P25RR   : in    std_logic;
    P25RO1  : out   std_logic;
    P25RO2  : out   std_logic;
    P25RO3  : out   std_logic;
    P25RO4  : out   std_logic;
    P25RO5  : out   std_logic;

    P26CI1  : in    std_logic;
    P26CL   : in    std_logic;
    P26CR   : in    std_logic;
    P26CO   : out   std_logic;
    P26CTI  : in    std_logic;
    P26CTO  : out   std_logic;
    P26EI1  : in    std_logic;
    P26EI2  : in    std_logic;
    P26EI3  : in    std_logic;
    P26EI4  : in    std_logic;
    P26EI5  : in    std_logic;
    P26EL   : in    std_logic;
    P26ER   : in    std_logic;
    P26EO   : out   std_logic;
    P26RI   : in    std_logic;
    P26RL   : in    std_logic;
    P26RR   : in    std_logic;
    P26RO1  : out   std_logic;
    P26RO2  : out   std_logic;
    P26RO3  : out   std_logic;
    P26RO4  : out   std_logic;
    P26RO5  : out   std_logic;

    P27CI1  : in    std_logic;
    P27CL   : in    std_logic;
    P27CR   : in    std_logic;
    P27CO   : out   std_logic;
    P27CTI  : in    std_logic;
    P27CTO  : out   std_logic;
    P27EI1  : in    std_logic;
    P27EI2  : in    std_logic;
    P27EI3  : in    std_logic;
    P27EI4  : in    std_logic;
    P27EI5  : in    std_logic;
    P27EL   : in    std_logic;
    P27ER   : in    std_logic;
    P27EO   : out   std_logic;
    P27RI   : in    std_logic;
    P27RL   : in    std_logic;
    P27RR   : in    std_logic;
    P27RO1  : out   std_logic;
    P27RO2  : out   std_logic;
    P27RO3  : out   std_logic;
    P27RO4  : out   std_logic;
    P27RO5  : out   std_logic;

    P28CI1  : in    std_logic;
    P28CL   : in    std_logic;
    P28CR   : in    std_logic;
    P28CO   : out   std_logic;
    P28CTI  : in    std_logic;
    P28CTO  : out   std_logic;
    P28EI1  : in    std_logic;
    P28EI2  : in    std_logic;
    P28EI3  : in    std_logic;
    P28EI4  : in    std_logic;
    P28EI5  : in    std_logic;
    P28EL   : in    std_logic;
    P28ER   : in    std_logic;
    P28EO   : out   std_logic;
    P28RI   : in    std_logic;
    P28RL   : in    std_logic;
    P28RR   : in    std_logic;
    P28RO1  : out   std_logic;
    P28RO2  : out   std_logic;
    P28RO3  : out   std_logic;
    P28RO4  : out   std_logic;
    P28RO5  : out   std_logic;

    P29CI1  : in    std_logic;
    P29CL   : in    std_logic;
    P29CR   : in    std_logic;
    P29CO   : out   std_logic;
    P29CTI  : in    std_logic;
    P29CTO  : out   std_logic;
    P29EI1  : in    std_logic;
    P29EI2  : in    std_logic;
    P29EI3  : in    std_logic;
    P29EI4  : in    std_logic;
    P29EI5  : in    std_logic;
    P29EL   : in    std_logic;
    P29ER   : in    std_logic;
    P29EO   : out   std_logic;
    P29RI   : in    std_logic;
    P29RL   : in    std_logic;
    P29RR   : in    std_logic;
    P29RO1  : out   std_logic;
    P29RO2  : out   std_logic;
    P29RO3  : out   std_logic;
    P29RO4  : out   std_logic;
    P29RO5  : out   std_logic;

    P30CI1  : in    std_logic;
    P30CL   : in    std_logic;
    P30CR   : in    std_logic;
    P30CO   : out   std_logic;
    P30CTI  : in    std_logic;
    P30CTO  : out   std_logic;
    P30EI1  : in    std_logic;
    P30EI2  : in    std_logic;
    P30EI3  : in    std_logic;
    P30EI4  : in    std_logic;
    P30EI5  : in    std_logic;
    P30EL   : in    std_logic;
    P30ER   : in    std_logic;
    P30EO   : out   std_logic;
    P30RI   : in    std_logic;
    P30RL   : in    std_logic;
    P30RR   : in    std_logic;
    P30RO1  : out   std_logic;
    P30RO2  : out   std_logic;
    P30RO3  : out   std_logic;
    P30RO4  : out   std_logic;
    P30RO5  : out   std_logic
);
end NX_IOM;

-- =================================================================================================
--   NX_IOM_CONTROL_M definition                                                         2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_CONTROL_M is
generic (
    mode_side1   : integer := 0;
    sel_clkw_rx1 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx1 : bit := '0';
    div_tx1      : bit_vector(3 downto 0) := "0000";
    div_rx1      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk1 : bit := '0';
    latency1     : bit := '0';
    mode_side2   : integer := 0;
    sel_clkw_rx2 : bit_vector(1 downto 0) := "00";
    sel_clkr_rx2 : bit := '0';
    div_tx2      : bit_vector(3 downto 0) := "0000";
    div_rx2      : bit_vector(3 downto 0) := "0000";
    inv_di_fclk2 : bit := '0';
    latency2     : bit := '0';
    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';
    mode_rpath   : string := "";
    mode_epath   : string := "";
    mode_cpath   : string := "";
    mode_tpath   : string := "";
    mode_io_cal  : bit    := '0';
    location  : string    := ""
);
port(
    RTCK1   : in    std_logic;
    RRCK1   : in    std_logic;
    WTCK1   : in    std_logic;
    WRCK1   : in    std_logic;
    RTCK2   : in    std_logic;
    RRCK2   : in    std_logic;
    WTCK2   : in    std_logic;
    WRCK2   : in    std_logic;
    CTCK    : in    std_logic;

    C1TW    : in    std_logic;
    C1TS    : in    std_logic;
    C1RW1   : in    std_logic;
    C1RW2   : in    std_logic;
    C1RW3   : in    std_logic;
    C1RNE   : in    std_logic;
    C1RS    : in    std_logic;
    C2TW    : in    std_logic;
    C2TS    : in    std_logic;
    C2RW1   : in    std_logic;
    C2RW2   : in    std_logic;
    C2RW3   : in    std_logic;
    C2RNE   : in    std_logic;
    C2RS    : in    std_logic;
    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;
    DC      : in    std_logic;
    CCK     : in    std_logic;
    DCK     : in    std_logic;
    DRI1    : in    std_logic;
    DRI2    : in    std_logic;
    DRI3    : in    std_logic;
    DRI4    : in    std_logic;
    DRI5    : in    std_logic;
    DRI6    : in    std_logic;
    DRA1    : in    std_logic;
    DRA2    : in    std_logic;
    DRA3    : in    std_logic;
    DRA4    : in    std_logic;
    DRA5    : in    std_logic;
    DRA6    : in    std_logic;
    DRL     : in    std_logic;
    DOS     : in    std_logic;
    DOG     : in    std_logic;
    DIS     : in    std_logic;
    DIG     : in    std_logic;
    DPAS    : in    std_logic;
    DPAG    : in    std_logic;
    DQSS    : in    std_logic;
    DQSG    : in    std_logic;
    DS1     : in    std_logic;
    DS2     : in    std_logic;
    CAD1    : in    std_logic;
    CAD2    : in    std_logic;
    CAD3    : in    std_logic;
    CAD4    : in    std_logic;
    CAD5    : in    std_logic;
    CAD6    : in    std_logic;
    CAP1    : in    std_logic;
    CAP2    : in    std_logic;
    CAP3    : in    std_logic;
    CAP4    : in    std_logic;
    CAN1    : in    std_logic;
    CAN2    : in    std_logic;
    CAN3    : in    std_logic;
    CAN4    : in    std_logic;
    CAT1    : in    std_logic;
    CAT2    : in    std_logic;
    CAT3    : in    std_logic;
    CAT4    : in    std_logic;
    SPI1    : in    std_logic;
    SPI2    : in    std_logic;
    SPI3    : in    std_logic;
    CKO1    : out   std_logic;
    CKO2    : out   std_logic;
    FLD     : out   std_logic;
    FLG     : out   std_logic;
    C1RED   : out   std_logic;
    C2RED   : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;
    CAL     : out   std_logic;

    LINK1  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK2  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK3  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK4  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK5  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK6  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK7  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK8  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK9  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK10 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK11 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK12 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK13 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK14 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK15 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK16 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK17 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK18 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK19 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK20 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK21 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK22 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK23 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK24 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK25 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK26 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK27 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK28 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK29 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK30 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK31 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK32 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK33 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK34 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_CONTROL_M;
-- =================================================================================================
--   NX_IOM_DRIVER_U definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_DRIVER_U is
generic (
    epath_edge      : bit := '0';
    epath_init      : bit := '0';
    epath_load      : bit := '0';
    epath_mode      : bit_vector(3 downto 0) := "0000";
    epath_sync      : bit := '0';
    epath_type      : bit := '0';
    epath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    rpath_edge      : bit := '0';
    rpath_init      : bit := '0';
    rpath_load      : bit := '0';
    rpath_mode      : bit_vector(3 downto 0) := "0000";
    rpath_sync      : bit := '0';
    rpath_type      : bit := '0';
    rpath_dynamic   : bit := '0'; --0: off/fixed delay, 1: dynamic delay

    cpath_edge      : bit := '0';
    cpath_init      : bit := '0';
    cpath_load      : bit := '0';
    cpath_mode      : bit_vector(3 downto 0) := "0000";
    cpath_sync      : bit := '0';
    cpath_type      : bit := '0';
    cpath_inv       : bit := '0';

    tpath_mode      : bit := '0';

    location        : string := "";
    chained         : bit    := '0';
    symbol          : string := ""
);
port (
    EI1  : in  std_logic;
    EI2  : in  std_logic;
    EI3  : in  std_logic;
    EI4  : in  std_logic;
    EI5  : in  std_logic;
    EI6  : in  std_logic;
    EI7  : in  std_logic;
    EI8  : in  std_logic;
    EL   : in  std_logic;
    ER   : in  std_logic;
    CI1  : in  std_logic;
    CL   : in  std_logic;
    CR   : in  std_logic;
    RI   : in  std_logic;
    RL   : in  std_logic;
    RR   : in  std_logic;
    CO   : out std_logic;
    CTI  : in  std_logic;
    CTO  : out std_logic;
    EO   : out std_logic;
    RO1  : out std_logic;
    RO2  : out std_logic;
    RO3  : out std_logic;
    RO4  : out std_logic;
    RO5  : out std_logic;
    RO6  : out std_logic;
    RO7  : out std_logic;
    RO8  : out std_logic;
    LINK : inout  std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_DRIVER_U;

-- =================================================================================================
--   NX_IOM_BIN2GRP definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_BIN2GRP is
port (
    LA    : in  std_logic_vector(5 downto 0);
    DS    : in  std_logic_vector(1 downto 0);

    GS    : in  std_logic;

    GVON  : out std_logic_vector(2 downto 0);
    GVIN  : out std_logic_vector(2 downto 0);
    GVDN  : out std_logic_vector(2 downto 0);
    PA    : out std_logic_vector(3 downto 0)
);
end NX_IOM_BIN2GRP;

architecture NX_RTL of NX_IOM_BIN2GRP is

    signal G    : std_logic_vector(2 downto 0);
    signal GSON : std_logic;
    signal GSIN : std_logic;
    signal GSDN : std_logic;

    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "LIB";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_BIN2GRP";

begin

GSON <= (not GS) when DS = "00" else '1';
GSIN <= (not GS) when DS = "01" else '1';
GSDN <= (not GS) when DS = "10" else '1';

process (LA)
begin
    case LA is

	when "000000" => PA <= "0001"; G <= "001";  -- Pad P01
	when "000001" => PA <= "0010"; G <= "001";  -- Pad P02
	when "000010" => PA <= "0011"; G <= "001";  -- Pad P03
	when "000011" => PA <= "0100"; G <= "001";  -- Pad P04
 
	when "000100" => PA <= "0101"; G <= "001";  -- Pad P05
	when "000101" => PA <= "0110"; G <= "001";  -- Pad P06
	when "000110" => PA <= "0111"; G <= "001";  -- Pad P07
	when "000111" => PA <= "1000"; G <= "001";  -- Pad P08

	when "001000" => PA <= "1001"; G <= "001";  -- Pad P09
	when "001001" => PA <= "1010"; G <= "001";  -- Pad P10
	when "001010" => PA <= "1011"; G <= "001";  -- Pad P11

--

	when "001011" => PA <= "0001"; G <= "001";  -- Pad P12
	when "001100" => PA <= "0010"; G <= "010";  -- Pad P13
	when "001101" => PA <= "0011"; G <= "010";  -- Pad P14
	when "001110" => PA <= "0100"; G <= "010";  -- Pad P15

	when "001111" => PA <= "0101"; G <= "010";  -- Pad P16
	when "010000" => PA <= "0110"; G <= "010";  -- Pad P17
	when "010001" => PA <= "0111"; G <= "010";  -- Pad P18
	when "010010" => PA <= "1000"; G <= "010";  -- Pad P19

	when "010011" => PA <= "1001"; G <= "010";  -- Pad P20
	when "010100" => PA <= "1010"; G <= "010";  -- Pad P21
	when "010101" => PA <= "1011"; G <= "010";  -- Pad P22

--

	when "010110" => PA <= "0001"; G <= "100";  -- Pad P23
	when "010111" => PA <= "0010"; G <= "100";  -- Pad P24
	when "011000" => PA <= "0011"; G <= "100";  -- Pad P25
	when "011001" => PA <= "0100"; G <= "100";  -- Pad P26

	when "011010" => PA <= "0101"; G <= "100";  -- Pad P27
	when "011011" => PA <= "0110"; G <= "100";  -- Pad P28
	when "011100" => PA <= "0111"; G <= "100";  -- Pad P29
	when "011101" => PA <= "1000"; G <= "100";  -- Pad P30

	when "011110" => PA <= "1001"; G <= "100";  -- Pad P31
	when "011111" => PA <= "1010"; G <= "100";  -- Pad P32
	when "100000" => PA <= "1011"; G <= "100";  -- Pad P33
	when "100001" => PA <= "1100"; G <= "100";  -- Pad P34

	when others   => PA <= "0000"; G <= "000";  -- Pad P34
    end case;
end process;

    GVON(0) <= GSON or (not G(0));
    GVON(1) <= GSON or (not G(1));
    GVON(2) <= GSON or (not G(2));

    GVIN(0) <= GSIN or (not G(0));
    GVIN(1) <= GSIN or (not G(1));
    GVIN(2) <= GSIN or (not G(2));

    GVDN(0) <= GSDN or (not G(0));
    GVDN(1) <= GSDN or (not G(1));
    GVDN(2) <= GSDN or (not G(2));

end NX_RTL;

-- =================================================================================================
--   NX_IOM_SERDES definition                                                             2018/10/15
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_SERDES_U is
generic (
    data_size : integer range 2 to 10 := 5;
    location  : string := ""
);
port (
    FCK   : in std_logic;
    SCK   : in std_logic;
    LDRN   : in std_logic;

    DRWDS  : in std_logic;
    DRWEN  : in std_logic;
    DRE    : in std_logic;
    DRON   : in std_logic_vector(2 downto 0);
    DRIN   : in std_logic_vector(2 downto 0);
    DRDN   : in std_logic_vector(2 downto 0);
    DRA    : in std_logic_vector(3 downto 0);
    DRI   : in std_logic_vector(5 downto 0);

    FA     : in std_logic_vector(5 downto 0);
    FZ    : in std_logic;

    ALD    : out std_logic;
    ALT    : out std_logic;

    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0);

    FLD   : out std_logic;
    FLG   : out std_logic;

    LINK   : inout std_logic_vector(IOM_LINK_SIZE-1 downto 0)
);
end NX_IOM_SERDES_U;
-- =================================================================================================
--   NX_IOM_U definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_U is
generic (
    mode_side1        : integer := 0;
    div1         : bit_vector(2 downto 0) := "000";
    mode_side2        : integer := 0;
    div2         : bit_vector(2 downto 0) := "000";
    mode_side3        : integer := 0;
    div3         : bit_vector(2 downto 0) := "000";

    div_swrx1    : bit_vector(2 downto 0) := "000";
    div_swrx2    : bit_vector(2 downto 0) := "000";

    sel_ld_fck1  : bit_vector(1 downto 0) := "00";
    sel_ld_fck2  : bit_vector(1 downto 0) := "00";
    sel_ld_fck3  : bit_vector(1 downto 0) := "00";
    sel_sw_fck1  : bit_vector(1 downto 0) := "00";
    sel_sw_fck2  : bit_vector(1 downto 0) := "00";

    sel_dc_clk   : bit_vector(1 downto 0) := "00";

    inv_ld_sck1  : bit := '0';
    inv_ld_sck2  : bit := '0';
    inv_ld_sck3  : bit := '0';

    link_ld_12   : bit := '0';
    link_ld_23   : bit := '0';

    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';

    use_dc       : bit := '0';
    cal_delay1   : string := "";
    cal_delay2   : string := "";

    pads_dict    : string := "";
    pads_path    : string := ""
);
port(
    ALCK1   : in    std_logic;
    ALCK2   : in    std_logic;
    ALCK3   : in    std_logic;
    LDSCK1  : in    std_logic;
    LDSCK2  : in    std_logic;
    LDSCK3  : in    std_logic;
--  LDFCK1  : in    std_logic;	-- CONFIG
--  LDFCK2  : in    std_logic;	-- CONFIG
--  LDFCK3  : in    std_logic;	-- CONFIG
--  SWTX1CK : in    std_logic;	-- CONFIG
--  SWTX2CK : in    std_logic;	-- CONFIG
    SWRX1CK : in    std_logic;
    SWRX2CK : in    std_logic;
    FCK1    : in    std_logic;
    FCK2    : in    std_logic;
    FDCK    : in    std_logic;
    CCK     : in    std_logic;

    DQ1CI1  : in    std_logic;
    DQ1CI2  : in    std_logic;
    DQ1CI3  : in    std_logic;
    DQ1CI4  : in    std_logic;
    DQ1CI5  : in    std_logic;
    DQ1CI6  : in    std_logic;
    DQ1CI7  : in    std_logic;
    DQ1CI8  : in    std_logic;
    DQ2CI1  : in    std_logic;
    DQ2CI2  : in    std_logic;
    DQ2CI3  : in    std_logic;
    DQ2CI4  : in    std_logic;
    DQ2CI5  : in    std_logic;
    DQ2CI6  : in    std_logic;
    DQ2CI7  : in    std_logic;
    DQ2CI8  : in    std_logic;
    DQ3CI1  : in    std_logic;
    DQ3CI2  : in    std_logic;
    DQ3CI3  : in    std_logic;
    DQ3CI4  : in    std_logic;
    DQ3CI5  : in    std_logic;
    DQ3CI6  : in    std_logic;
    DQ3CI7  : in    std_logic;
    DQ3CI8  : in    std_logic;
    DQS1CI1 : in    std_logic;
    DQS1CI2 : in    std_logic;
    DQS1CI3 : in    std_logic;
    DQS1CI4 : in    std_logic;
    DQS1CI5 : in    std_logic;
    DQS1CI6 : in    std_logic;
    DQS1CI7 : in    std_logic;
    DQS1CI8 : in    std_logic;
    DQS2CI1 : in    std_logic;
    DQS2CI2 : in    std_logic;
    DQS2CI3 : in    std_logic;
    DQS2CI4 : in    std_logic;
    DQS2CI5 : in    std_logic;
    DQS2CI6 : in    std_logic;
    DQS2CI7 : in    std_logic;
    DQS2CI8 : in    std_logic;
    DQS3CI1 : in    std_logic;
    DQS3CI2 : in    std_logic;
    DQS3CI3 : in    std_logic;
    DQS3CI4 : in    std_logic;
    DQS3CI5 : in    std_logic;
    DQS3CI6 : in    std_logic;
    DQS3CI7 : in    std_logic;
    DQS3CI8 : in    std_logic;

    LD1RN   : in    std_logic;
    LD2RN   : in    std_logic;
    LD3RN   : in    std_logic;

    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;

    DCRN    : in    std_logic;
    LE      : in    std_logic;
    SE      : in    std_logic;

    DRI1     : in    std_logic;
    DRI2     : in    std_logic;
    DRI3     : in    std_logic;
    DRI4     : in    std_logic;
    DRI5     : in    std_logic;
    DRI6     : in    std_logic;
    DRA1     : in    std_logic;
    DRA2     : in    std_logic;
    DRA3     : in    std_logic;
    DRA4     : in    std_logic;

    DRO1CSN   : in    std_logic;
    DRO2CSN   : in    std_logic;
    DRO3CSN   : in    std_logic;
    DRI1CSN   : in    std_logic;
    DRI2CSN   : in    std_logic;
    DRI3CSN   : in    std_logic;
    DRDPA1CSN : in    std_logic;
    DRDPA2CSN : in    std_logic;
    DRDPA3CSN : in    std_logic;
    DRCCSN    : in    std_logic;
    DRWDS     : in    std_logic;
    DRWEN     : in    std_logic;
    DRE       : in    std_logic;

    CA1P1   : in    std_logic;
    CA1P2   : in    std_logic;
    CA1P3   : in    std_logic;
    CA1P4   : in    std_logic;
    CA2P1   : in    std_logic;
    CA2P2   : in    std_logic;
    CA2P3   : in    std_logic;
    CA2P4   : in    std_logic;
    CA1N1   : in    std_logic;
    CA1N2   : in    std_logic;
    CA1N3   : in    std_logic;
    CA1N4   : in    std_logic;
    CA2N1   : in    std_logic;
    CA2N2   : in    std_logic;
    CA2N3   : in    std_logic;
    CA2N4   : in    std_logic;
    CA1T1   : in    std_logic;
    CA1T2   : in    std_logic;
    CA1T3   : in    std_logic;
    CA1T4   : in    std_logic;
    CA2T1   : in    std_logic;
    CA2T2   : in    std_logic;
    CA2T3   : in    std_logic;
    CA2T4   : in    std_logic;
    CA1D1   : in    std_logic;
    CA1D2   : in    std_logic;
    CA1D3   : in    std_logic;
    CA1D4   : in    std_logic;
    CA1D5   : in    std_logic;
    CA1D6   : in    std_logic;
    CA2D1   : in    std_logic;
    CA2D2   : in    std_logic;
    CA2D3   : in    std_logic;
    CA2D4   : in    std_logic;
    CA2D5   : in    std_logic;
    CA2D6   : in    std_logic;

    CKO1    : out   std_logic;
    CKO2    : out   std_logic;

    FLD     : out   std_logic;
    FLG     : out   std_logic;
    AL1D    : out   std_logic;
    AL2D    : out   std_logic;
    AL3D    : out   std_logic;
    AL1T    : out   std_logic;
    AL2T    : out   std_logic;
    AL3T    : out   std_logic;
    DCL     : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;

    P1CI1   : in    std_logic;
    P1CL    : in    std_logic;
    P1CR    : in    std_logic;
    P1CO    : out   std_logic;
    P1CTI   : in    std_logic;
    P1CTO   : out   std_logic;
    P1EI1   : in    std_logic;
    P1EI2   : in    std_logic;
    P1EI3   : in    std_logic;
    P1EI4   : in    std_logic;
    P1EI5   : in    std_logic;
    P1EI6   : in    std_logic;
    P1EI7   : in    std_logic;
    P1EI8   : in    std_logic;

    P1EL    : in    std_logic;
    P1ER    : in    std_logic;
    P1EO    : out   std_logic;
    P1RI    : in    std_logic;
    P1RL    : in    std_logic;
    P1RR    : in    std_logic;
    P1RO1   : out   std_logic;
    P1RO2   : out   std_logic;
    P1RO3   : out   std_logic;
    P1RO4   : out   std_logic;
    P1RO5   : out   std_logic;
    P1RO6   : out   std_logic;
    P1RO7   : out   std_logic;
    P1RO8   : out   std_logic;

    P2CI1   : in    std_logic;
    P2CL    : in    std_logic;
    P2CR    : in    std_logic;
    P2CO    : out   std_logic;
    P2CTI   : in    std_logic;
    P2CTO   : out   std_logic;
    P2EI1   : in    std_logic;
    P2EI2   : in    std_logic;
    P2EI3   : in    std_logic;
    P2EI4   : in    std_logic;
    P2EI5   : in    std_logic;
    P2EI6   : in    std_logic;
    P2EI7   : in    std_logic;
    P2EI8   : in    std_logic;

    P2EL    : in    std_logic;
    P2ER    : in    std_logic;
    P2EO    : out   std_logic;
    P2RI    : in    std_logic;
    P2RL    : in    std_logic;
    P2RR    : in    std_logic;
    P2RO1   : out   std_logic;
    P2RO2   : out   std_logic;
    P2RO3   : out   std_logic;
    P2RO4   : out   std_logic;
    P2RO5   : out   std_logic;
    P2RO6   : out   std_logic;
    P2RO7   : out   std_logic;
    P2RO8   : out   std_logic;

    P3CI1   : in    std_logic;
    P3CL    : in    std_logic;
    P3CR    : in    std_logic;
    P3CO    : out   std_logic;
    P3CTI   : in    std_logic;
    P3CTO   : out   std_logic;
    P3EI1   : in    std_logic;
    P3EI2   : in    std_logic;
    P3EI3   : in    std_logic;
    P3EI4   : in    std_logic;
    P3EI5   : in    std_logic;
    P3EI6   : in    std_logic;
    P3EI7   : in    std_logic;
    P3EI8   : in    std_logic;

    P3EL    : in    std_logic;
    P3ER    : in    std_logic;
    P3EO    : out   std_logic;
    P3RI    : in    std_logic;
    P3RL    : in    std_logic;
    P3RR    : in    std_logic;
    P3RO1   : out   std_logic;
    P3RO2   : out   std_logic;
    P3RO3   : out   std_logic;
    P3RO4   : out   std_logic;
    P3RO5   : out   std_logic;
    P3RO6   : out   std_logic;
    P3RO7   : out   std_logic;
    P3RO8   : out   std_logic;

    P4CI1   : in    std_logic;
    P4CL    : in    std_logic;
    P4CR    : in    std_logic;
    P4CO    : out   std_logic;
    P4CTI   : in    std_logic;
    P4CTO   : out   std_logic;
    P4EI1   : in    std_logic;
    P4EI2   : in    std_logic;
    P4EI3   : in    std_logic;
    P4EI4   : in    std_logic;
    P4EI5   : in    std_logic;
    P4EI6   : in    std_logic;
    P4EI7   : in    std_logic;
    P4EI8   : in    std_logic;

    P4EL    : in    std_logic;
    P4ER    : in    std_logic;
    P4EO    : out   std_logic;
    P4RI    : in    std_logic;
    P4RL    : in    std_logic;
    P4RR    : in    std_logic;
    P4RO1   : out   std_logic;
    P4RO2   : out   std_logic;
    P4RO3   : out   std_logic;
    P4RO4   : out   std_logic;
    P4RO5   : out   std_logic;
    P4RO6   : out   std_logic;
    P4RO7   : out   std_logic;
    P4RO8   : out   std_logic;

    P5CI1   : in    std_logic;
    P5CL    : in    std_logic;
    P5CR    : in    std_logic;
    P5CO    : out   std_logic;
    P5CTI   : in    std_logic;
    P5CTO   : out   std_logic;
    P5EI1   : in    std_logic;
    P5EI2   : in    std_logic;
    P5EI3   : in    std_logic;
    P5EI4   : in    std_logic;
    P5EI5   : in    std_logic;
    P5EI6   : in    std_logic;
    P5EI7   : in    std_logic;
    P5EI8   : in    std_logic;

    P5EL    : in    std_logic;
    P5ER    : in    std_logic;
    P5EO    : out   std_logic;
    P5RI    : in    std_logic;
    P5RL    : in    std_logic;
    P5RR    : in    std_logic;
    P5RO1   : out   std_logic;
    P5RO2   : out   std_logic;
    P5RO3   : out   std_logic;
    P5RO4   : out   std_logic;
    P5RO5   : out   std_logic;
    P5RO6   : out   std_logic;
    P5RO7   : out   std_logic;
    P5RO8   : out   std_logic;

    P6CI1   : in    std_logic;
    P6CL    : in    std_logic;
    P6CR    : in    std_logic;
    P6CO    : out   std_logic;
    P6CTI   : in    std_logic;
    P6CTO   : out   std_logic;
    P6EI1   : in    std_logic;
    P6EI2   : in    std_logic;
    P6EI3   : in    std_logic;
    P6EI4   : in    std_logic;
    P6EI5   : in    std_logic;
    P6EI6   : in    std_logic;
    P6EI7   : in    std_logic;
    P6EI8   : in    std_logic;

    P6EL    : in    std_logic;
    P6ER    : in    std_logic;
    P6EO    : out   std_logic;
    P6RI    : in    std_logic;
    P6RL    : in    std_logic;
    P6RR    : in    std_logic;
    P6RO1   : out   std_logic;
    P6RO2   : out   std_logic;
    P6RO3   : out   std_logic;
    P6RO4   : out   std_logic;
    P6RO5   : out   std_logic;
    P6RO6   : out   std_logic;
    P6RO7   : out   std_logic;
    P6RO8   : out   std_logic;

    P7CI1   : in    std_logic;
    P7CL    : in    std_logic;
    P7CR    : in    std_logic;
    P7CO    : out   std_logic;
    P7CTI   : in    std_logic;
    P7CTO   : out   std_logic;
    P7EI1   : in    std_logic;
    P7EI2   : in    std_logic;
    P7EI3   : in    std_logic;
    P7EI4   : in    std_logic;
    P7EI5   : in    std_logic;
    P7EI6   : in    std_logic;
    P7EI7   : in    std_logic;
    P7EI8   : in    std_logic;

    P7EL    : in    std_logic;
    P7ER    : in    std_logic;
    P7EO    : out   std_logic;
    P7RI    : in    std_logic;
    P7RL    : in    std_logic;
    P7RR    : in    std_logic;
    P7RO1   : out   std_logic;
    P7RO2   : out   std_logic;
    P7RO3   : out   std_logic;
    P7RO4   : out   std_logic;
    P7RO5   : out   std_logic;
    P7RO6   : out   std_logic;
    P7RO7   : out   std_logic;
    P7RO8   : out   std_logic;

    P8CI1   : in    std_logic;
    P8CL    : in    std_logic;
    P8CR    : in    std_logic;
    P8CO    : out   std_logic;
    P8CTI   : in    std_logic;
    P8CTO   : out   std_logic;
    P8EI1   : in    std_logic;
    P8EI2   : in    std_logic;
    P8EI3   : in    std_logic;
    P8EI4   : in    std_logic;
    P8EI5   : in    std_logic;
    P8EI6   : in    std_logic;
    P8EI7   : in    std_logic;
    P8EI8   : in    std_logic;

    P8EL    : in    std_logic;
    P8ER    : in    std_logic;
    P8EO    : out   std_logic;
    P8RI    : in    std_logic;
    P8RL    : in    std_logic;
    P8RR    : in    std_logic;
    P8RO1   : out   std_logic;
    P8RO2   : out   std_logic;
    P8RO3   : out   std_logic;
    P8RO4   : out   std_logic;
    P8RO5   : out   std_logic;
    P8RO6   : out   std_logic;
    P8RO7   : out   std_logic;
    P8RO8   : out   std_logic;

    P9CI1   : in    std_logic;
    P9CL    : in    std_logic;
    P9CR    : in    std_logic;
    P9CO    : out   std_logic;
    P9CTI   : in    std_logic;
    P9CTO   : out   std_logic;
    P9EI1   : in    std_logic;
    P9EI2   : in    std_logic;
    P9EI3   : in    std_logic;
    P9EI4   : in    std_logic;
    P9EI5   : in    std_logic;
    P9EI6   : in    std_logic;
    P9EI7   : in    std_logic;
    P9EI8   : in    std_logic;

    P9EL    : in    std_logic;
    P9ER    : in    std_logic;
    P9EO    : out   std_logic;
    P9RI    : in    std_logic;
    P9RL    : in    std_logic;
    P9RR    : in    std_logic;
    P9RO1   : out   std_logic;
    P9RO2   : out   std_logic;
    P9RO3   : out   std_logic;
    P9RO4   : out   std_logic;
    P9RO5   : out   std_logic;
    P9RO6   : out   std_logic;
    P9RO7   : out   std_logic;
    P9RO8   : out   std_logic;

    P10CI1  : in    std_logic;
    P10CL   : in    std_logic;
    P10CR   : in    std_logic;
    P10CO   : out   std_logic;
    P10CTI  : in    std_logic;
    P10CTO  : out   std_logic;
    P10EI1  : in    std_logic;
    P10EI2  : in    std_logic;
    P10EI3  : in    std_logic;
    P10EI4  : in    std_logic;
    P10EI5  : in    std_logic;
    P10EI6  : in    std_logic;
    P10EI7  : in    std_logic;
    P10EI8  : in    std_logic;

    P10EL   : in    std_logic;
    P10ER   : in    std_logic;
    P10EO   : out   std_logic;
    P10RI   : in    std_logic;
    P10RL   : in    std_logic;
    P10RR   : in    std_logic;
    P10RO1  : out   std_logic;
    P10RO2  : out   std_logic;
    P10RO3  : out   std_logic;
    P10RO4  : out   std_logic;
    P10RO5  : out   std_logic;
    P10RO6  : out   std_logic;
    P10RO7  : out   std_logic;
    P10RO8  : out   std_logic;

    P11CI1  : in    std_logic;
    
    P11CL   : in    std_logic;
    P11CR   : in    std_logic;
    P11CO   : out   std_logic;
    P11CTI  : in    std_logic;
    P11CTO  : out   std_logic;
    P11EI1  : in    std_logic;
    P11EI2  : in    std_logic;
    P11EI3  : in    std_logic;
    P11EI4  : in    std_logic;
    P11EI5  : in    std_logic;
    P11EI6  : in    std_logic;
    P11EI7  : in    std_logic;
    P11EI8  : in    std_logic;

    P11EL   : in    std_logic;
    P11ER   : in    std_logic;
    P11EO   : out   std_logic;
    P11RI   : in    std_logic;
    P11RL   : in    std_logic;
    P11RR   : in    std_logic;
    P11RO1  : out   std_logic;
    P11RO2  : out   std_logic;
    P11RO3  : out   std_logic;
    P11RO4  : out   std_logic;
    P11RO5  : out   std_logic;
    P11RO6  : out   std_logic;
    P11RO7  : out   std_logic;
    P11RO8  : out   std_logic;

    P12CI1  : in    std_logic;
    P12CL   : in    std_logic;
    P12CR   : in    std_logic;
    P12CO   : out   std_logic;
    P12CTI  : in    std_logic;
    P12CTO  : out   std_logic;
    P12EI1  : in    std_logic;
    P12EI2  : in    std_logic;
    P12EI3  : in    std_logic;
    P12EI4  : in    std_logic;
    P12EI5  : in    std_logic;
    P12EI6  : in    std_logic;
    P12EI7  : in    std_logic;
    P12EI8  : in    std_logic;

    P12EL   : in    std_logic;
    P12ER   : in    std_logic;
    P12EO   : out   std_logic;
    P12RI   : in    std_logic;
    P12RL   : in    std_logic;
    P12RR   : in    std_logic;
    P12RO1  : out   std_logic;
    P12RO2  : out   std_logic;
    P12RO3  : out   std_logic;
    P12RO4  : out   std_logic;
    P12RO5  : out   std_logic;
    P12RO6  : out   std_logic;
    P12RO7  : out   std_logic;
    P12RO8  : out   std_logic;

    P13CI1  : in    std_logic;
    P13CL   : in    std_logic;
    P13CR   : in    std_logic;
    P13CO   : out   std_logic;
    P13CTI  : in    std_logic;
    P13CTO  : out   std_logic;
    P13EI1  : in    std_logic;
    P13EI2  : in    std_logic;
    P13EI3  : in    std_logic;
    P13EI4  : in    std_logic;
    P13EI5  : in    std_logic;
    P13EI6  : in    std_logic;
    P13EI7  : in    std_logic;
    P13EI8  : in    std_logic;

    P13EL   : in    std_logic;
    P13ER   : in    std_logic;
    P13EO   : out   std_logic;
    P13RI   : in    std_logic;
    P13RL   : in    std_logic;
    P13RR   : in    std_logic;
    P13RO1  : out   std_logic;
    P13RO2  : out   std_logic;
    P13RO3  : out   std_logic;
    P13RO4  : out   std_logic;
    P13RO5  : out   std_logic;
    P13RO6  : out   std_logic;
    P13RO7  : out   std_logic;
    P13RO8  : out   std_logic;

    P14CI1  : in    std_logic;
    P14CL   : in    std_logic;
    P14CR   : in    std_logic;
    P14CO   : out   std_logic;
    P14CTI  : in    std_logic;
    P14CTO  : out   std_logic;
    P14EI1  : in    std_logic;
    P14EI2  : in    std_logic;
    P14EI3  : in    std_logic;
    P14EI4  : in    std_logic;
    P14EI5  : in    std_logic;
    P14EI6  : in    std_logic;
    P14EI7  : in    std_logic;
    P14EI8  : in    std_logic;

    P14EL   : in    std_logic;
    P14ER   : in    std_logic;
    P14EO   : out   std_logic;
    P14RI   : in    std_logic;
    P14RL   : in    std_logic;
    P14RR   : in    std_logic;
    P14RO1  : out   std_logic;
    P14RO2  : out   std_logic;
    P14RO3  : out   std_logic;
    P14RO4  : out   std_logic;
    P14RO5  : out   std_logic;
    P14RO6  : out   std_logic;
    P14RO7  : out   std_logic;
    P14RO8  : out   std_logic;

    P15CI1  : in    std_logic;
    P15CL   : in    std_logic;
    P15CR   : in    std_logic;
    P15CO   : out   std_logic;
    P15CTI  : in    std_logic;
    P15CTO  : out   std_logic;
    P15EI1  : in    std_logic;
    P15EI2  : in    std_logic;
    P15EI3  : in    std_logic;
    P15EI4  : in    std_logic;
    P15EI5  : in    std_logic;
    P15EI6  : in    std_logic;
    P15EI7  : in    std_logic;
    P15EI8  : in    std_logic;

    P15EL   : in    std_logic;
    P15ER   : in    std_logic;
    P15EO   : out   std_logic;
    P15RI   : in    std_logic;
    P15RL   : in    std_logic;
    P15RR   : in    std_logic;
    P15RO1  : out   std_logic;
    P15RO2  : out   std_logic;
    P15RO3  : out   std_logic;
    P15RO4  : out   std_logic;
    P15RO5  : out   std_logic;
    P15RO6  : out   std_logic;
    P15RO7  : out   std_logic;
    P15RO8  : out   std_logic;

    P16CI1  : in    std_logic;
    P16CL   : in    std_logic;
    P16CR   : in    std_logic;
    P16CO   : out   std_logic;
    P16CTI  : in    std_logic;
    P16CTO  : out   std_logic;
    P16EI1  : in    std_logic;
    P16EI2  : in    std_logic;
    P16EI3  : in    std_logic;
    P16EI4  : in    std_logic;
    P16EI5  : in    std_logic;
    P16EI6  : in    std_logic;
    P16EI7  : in    std_logic;
    P16EI8  : in    std_logic;

    P16EL   : in    std_logic;
    P16ER   : in    std_logic;
    P16EO   : out   std_logic;
    P16RI   : in    std_logic;
    P16RL   : in    std_logic;
    P16RR   : in    std_logic;
    P16RO1  : out   std_logic;
    P16RO2  : out   std_logic;
    P16RO3  : out   std_logic;
    P16RO4  : out   std_logic;
    P16RO5  : out   std_logic;
    P16RO6  : out   std_logic;
    P16RO7  : out   std_logic;
    P16RO8  : out   std_logic;

    P17CI1  : in    std_logic;
    P17CL   : in    std_logic;
    P17CR   : in    std_logic;
    P17CO   : out   std_logic;
    P17CTI  : in    std_logic;
    P17CTO  : out   std_logic;
    P17EI1  : in    std_logic;
    P17EI2  : in    std_logic;
    P17EI3  : in    std_logic;
    P17EI4  : in    std_logic;
    P17EI5  : in    std_logic;
    P17EI6  : in    std_logic;
    P17EI7  : in    std_logic;
    P17EI8  : in    std_logic;

    P17EL   : in    std_logic;
    P17ER   : in    std_logic;
    P17EO   : out   std_logic;
    P17RI   : in    std_logic;
    P17RL   : in    std_logic;
    P17RR   : in    std_logic;
    P17RO1  : out   std_logic;
    P17RO2  : out   std_logic;
    P17RO3  : out   std_logic;
    P17RO4  : out   std_logic;
    P17RO5  : out   std_logic;
    P17RO6  : out   std_logic;
    P17RO7  : out   std_logic;
    P17RO8  : out   std_logic;

    P18CI1  : in    std_logic;
    P18CL   : in    std_logic;
    P18CR   : in    std_logic;
    P18CO   : out   std_logic;
    P18CTI  : in    std_logic;
    P18CTO  : out   std_logic;
    P18EI1  : in    std_logic;
    P18EI2  : in    std_logic;
    P18EI3  : in    std_logic;
    P18EI4  : in    std_logic;
    P18EI5  : in    std_logic;
    P18EI6  : in    std_logic;
    P18EI7  : in    std_logic;
    P18EI8  : in    std_logic;

    P18EL   : in    std_logic;
    P18ER   : in    std_logic;
    P18EO   : out   std_logic;
    P18RI   : in    std_logic;
    P18RL   : in    std_logic;
    P18RR   : in    std_logic;
    P18RO1  : out   std_logic;
    P18RO2  : out   std_logic;
    P18RO3  : out   std_logic;
    P18RO4  : out   std_logic;
    P18RO5  : out   std_logic;
    P18RO6  : out   std_logic;
    P18RO7  : out   std_logic;
    P18RO8  : out   std_logic;

    P19CI1  : in    std_logic;
    P19CL   : in    std_logic;
    P19CR   : in    std_logic;
    P19CO   : out   std_logic;
    P19CTI  : in    std_logic;
    P19CTO  : out   std_logic;
    P19EI1  : in    std_logic;
    P19EI2  : in    std_logic;
    P19EI3  : in    std_logic;
    P19EI4  : in    std_logic;
    P19EI5  : in    std_logic;
    P19EI6  : in    std_logic;
    P19EI7  : in    std_logic;
    P19EI8  : in    std_logic;

    P19EL   : in    std_logic;
    P19ER   : in    std_logic;
    P19EO   : out   std_logic;
    P19RI   : in    std_logic;
    P19RL   : in    std_logic;
    P19RR   : in    std_logic;
    P19RO1  : out   std_logic;
    P19RO2  : out   std_logic;
    P19RO3  : out   std_logic;
    P19RO4  : out   std_logic;
    P19RO5  : out   std_logic;
    P19RO6  : out   std_logic;
    P19RO7  : out   std_logic;
    P19RO8  : out   std_logic;

    P20CI1  : in    std_logic;
    P20CL   : in    std_logic;
    P20CR   : in    std_logic;
    P20CO   : out   std_logic;
    P20CTI  : in    std_logic;
    P20CTO  : out   std_logic;
    P20EI1  : in    std_logic;
    P20EI2  : in    std_logic;
    P20EI3  : in    std_logic;
    P20EI4  : in    std_logic;
    P20EI5  : in    std_logic;
    P20EI6  : in    std_logic;
    P20EI7  : in    std_logic;
    P20EI8  : in    std_logic;

    P20EL   : in    std_logic;
    P20ER   : in    std_logic;
    P20EO   : out   std_logic;
    P20RI   : in    std_logic;
    P20RL   : in    std_logic;
    P20RR   : in    std_logic;
    P20RO1  : out   std_logic;
    P20RO2  : out   std_logic;
    P20RO3  : out   std_logic;
    P20RO4  : out   std_logic;
    P20RO5  : out   std_logic;
    P20RO6  : out   std_logic;
    P20RO7  : out   std_logic;
    P20RO8  : out   std_logic;

    P21CI1  : in    std_logic;
    P21CL   : in    std_logic;
    P21CR   : in    std_logic;
    P21CO   : out   std_logic;
    P21CTI  : in    std_logic;
    P21CTO  : out   std_logic;
    P21EI1  : in    std_logic;
    P21EI2  : in    std_logic;
    P21EI3  : in    std_logic;
    P21EI4  : in    std_logic;
    P21EI5  : in    std_logic;
    P21EI6  : in    std_logic;
    P21EI7  : in    std_logic;
    P21EI8  : in    std_logic;

    P21EL   : in    std_logic;
    P21ER   : in    std_logic;
    P21EO   : out   std_logic;
    P21RI   : in    std_logic;
    P21RL   : in    std_logic;
    P21RR   : in    std_logic;
    P21RO1  : out   std_logic;
    P21RO2  : out   std_logic;
    P21RO3  : out   std_logic;
    P21RO4  : out   std_logic;
    P21RO5  : out   std_logic;
    P21RO6  : out   std_logic;
    P21RO7  : out   std_logic;
    P21RO8  : out   std_logic;

    P22CI1  : in    std_logic;
    P22CL   : in    std_logic;
    P22CR   : in    std_logic;
    P22CO   : out   std_logic;
    P22CTI  : in    std_logic;
    P22CTO  : out   std_logic;
    P22EI1  : in    std_logic;
    P22EI2  : in    std_logic;
    P22EI3  : in    std_logic;
    P22EI4  : in    std_logic;
    P22EI5  : in    std_logic;
    P22EI6  : in    std_logic;
    P22EI7  : in    std_logic;
    P22EI8  : in    std_logic;

    P22EL   : in    std_logic;
    P22ER   : in    std_logic;
    P22EO   : out   std_logic;
    P22RI   : in    std_logic;
    P22RL   : in    std_logic;
    P22RR   : in    std_logic;
    P22RO1  : out   std_logic;
    P22RO2  : out   std_logic;
    P22RO3  : out   std_logic;
    P22RO4  : out   std_logic;
    P22RO5  : out   std_logic;
    P22RO6  : out   std_logic;
    P22RO7  : out   std_logic;
    P22RO8  : out   std_logic;

    P23CI1  : in    std_logic;
    P23CL   : in    std_logic;
    P23CR   : in    std_logic;
    P23CO   : out   std_logic;
    P23CTI  : in    std_logic;
    P23CTO  : out   std_logic;
    P23EI1  : in    std_logic;
    P23EI2  : in    std_logic;
    P23EI3  : in    std_logic;
    P23EI4  : in    std_logic;
    P23EI5  : in    std_logic;
    P23EI6  : in    std_logic;
    P23EI7  : in    std_logic;
    P23EI8  : in    std_logic;

    P23EL   : in    std_logic;
    P23ER   : in    std_logic;
    P23EO   : out   std_logic;
    P23RI   : in    std_logic;
    P23RL   : in    std_logic;
    P23RR   : in    std_logic;
    P23RO1  : out   std_logic;
    P23RO2  : out   std_logic;
    P23RO3  : out   std_logic;
    P23RO4  : out   std_logic;
    P23RO5  : out   std_logic;
    P23RO6  : out   std_logic;
    P23RO7  : out   std_logic;
    P23RO8  : out   std_logic;

    P24CI1  : in    std_logic;
    P24CL   : in    std_logic;
    P24CR   : in    std_logic;
    P24CO   : out   std_logic;
    P24CTI  : in    std_logic;
    P24CTO  : out   std_logic;
    P24EI1  : in    std_logic;
    P24EI2  : in    std_logic;
    P24EI3  : in    std_logic;
    P24EI4  : in    std_logic;
    P24EI5  : in    std_logic;
    P24EI6  : in    std_logic;
    P24EI7  : in    std_logic;
    P24EI8  : in    std_logic;

    P24EL   : in    std_logic;
    P24ER   : in    std_logic;
    P24EO   : out   std_logic;
    P24RI   : in    std_logic;
    P24RL   : in    std_logic;
    P24RR   : in    std_logic;
    P24RO1  : out   std_logic;
    P24RO2  : out   std_logic;
    P24RO3  : out   std_logic;
    P24RO4  : out   std_logic;
    P24RO5  : out   std_logic;
    P24RO6  : out   std_logic;
    P24RO7  : out   std_logic;
    P24RO8  : out   std_logic;

    P25CI1  : in    std_logic;
    P25CL   : in    std_logic;
    P25CR   : in    std_logic;
    P25CO   : out   std_logic;
    P25CTI  : in    std_logic;
    P25CTO  : out   std_logic;
    P25EI1  : in    std_logic;
    P25EI2  : in    std_logic;
    P25EI3  : in    std_logic;
    P25EI4  : in    std_logic;
    P25EI5  : in    std_logic;
    P25EI6  : in    std_logic;
    P25EI7  : in    std_logic;
    P25EI8  : in    std_logic;

    P25EL   : in    std_logic;
    P25ER   : in    std_logic;
    P25EO   : out   std_logic;
    P25RI   : in    std_logic;
    P25RL   : in    std_logic;
    P25RR   : in    std_logic;
    P25RO1  : out   std_logic;
    P25RO2  : out   std_logic;
    P25RO3  : out   std_logic;
    P25RO4  : out   std_logic;
    P25RO5  : out   std_logic;
    P25RO6  : out   std_logic;
    P25RO7  : out   std_logic;
    P25RO8  : out   std_logic;

    P26CI1  : in    std_logic;
    P26CL   : in    std_logic;
    P26CR   : in    std_logic;
    P26CO   : out   std_logic;
    P26CTI  : in    std_logic;
    P26CTO  : out   std_logic;
    P26EI1  : in    std_logic;
    P26EI2  : in    std_logic;
    P26EI3  : in    std_logic;
    P26EI4  : in    std_logic;
    P26EI5  : in    std_logic;
    P26EI6  : in    std_logic;
    P26EI7  : in    std_logic;
    P26EI8  : in    std_logic;

    P26EL   : in    std_logic;
    P26ER   : in    std_logic;
    P26EO   : out   std_logic;
    P26RI   : in    std_logic;
    P26RL   : in    std_logic;
    P26RR   : in    std_logic;
    P26RO1  : out   std_logic;
    P26RO2  : out   std_logic;
    P26RO3  : out   std_logic;
    P26RO4  : out   std_logic;
    P26RO5  : out   std_logic;
    P26RO6  : out   std_logic;
    P26RO7  : out   std_logic;
    P26RO8  : out   std_logic;

    P27CI1  : in    std_logic;
    P27CL   : in    std_logic;
    P27CR   : in    std_logic;
    P27CO   : out   std_logic;
    P27CTI  : in    std_logic;
    P27CTO  : out   std_logic;
    P27EI1  : in    std_logic;
    P27EI2  : in    std_logic;
    P27EI3  : in    std_logic;
    P27EI4  : in    std_logic;
    P27EI5  : in    std_logic;
    P27EI6  : in    std_logic;
    P27EI7  : in    std_logic;
    P27EI8  : in    std_logic;

    P27EL   : in    std_logic;
    P27ER   : in    std_logic;
    P27EO   : out   std_logic;
    P27RI   : in    std_logic;
    P27RL   : in    std_logic;
    P27RR   : in    std_logic;
    P27RO1  : out   std_logic;
    P27RO2  : out   std_logic;
    P27RO3  : out   std_logic;
    P27RO4  : out   std_logic;
    P27RO5  : out   std_logic;
    P27RO6  : out   std_logic;
    P27RO7  : out   std_logic;
    P27RO8  : out   std_logic;

    P28CI1  : in    std_logic;
    P28CL   : in    std_logic;
    P28CR   : in    std_logic;
    P28CO   : out   std_logic;
    P28CTI  : in    std_logic;
    P28CTO  : out   std_logic;
    P28EI1  : in    std_logic;
    P28EI2  : in    std_logic;
    P28EI3  : in    std_logic;
    P28EI4  : in    std_logic;
    P28EI5  : in    std_logic;
    P28EI6  : in    std_logic;
    P28EI7  : in    std_logic;
    P28EI8  : in    std_logic;
    P28EL   : in    std_logic;
    P28ER   : in    std_logic;
    P28EO   : out   std_logic;
    P28RI   : in    std_logic;
    P28RL   : in    std_logic;
    P28RR   : in    std_logic;
    P28RO1  : out   std_logic;
    P28RO2  : out   std_logic;
    P28RO3  : out   std_logic;
    P28RO4  : out   std_logic;
    P28RO5  : out   std_logic;
    P28RO6  : out   std_logic;
    P28RO7  : out   std_logic;
    P28RO8  : out   std_logic;

    P29CI1  : in    std_logic;
    P29CL   : in    std_logic;
    P29CR   : in    std_logic;
    P29CO   : out   std_logic;
    P29CTI  : in    std_logic;
    P29CTO  : out   std_logic;
    P29EI1  : in    std_logic;
    P29EI2  : in    std_logic;
    P29EI3  : in    std_logic;
    P29EI4  : in    std_logic;
    P29EI5  : in    std_logic;
    P29EI6  : in    std_logic;
    P29EI7  : in    std_logic;
    P29EI8  : in    std_logic;
    P29EL   : in    std_logic;
    P29ER   : in    std_logic;
    P29EO   : out   std_logic;
    P29RI   : in    std_logic;
    P29RL   : in    std_logic;
    P29RR   : in    std_logic;
    P29RO1  : out   std_logic;
    P29RO2  : out   std_logic;
    P29RO3  : out   std_logic;
    P29RO4  : out   std_logic;
    P29RO5  : out   std_logic;
    P29RO6  : out   std_logic;
    P29RO7  : out   std_logic;
    P29RO8  : out   std_logic;

    P30CI1  : in    std_logic;
    P30CL   : in    std_logic;
    P30CR   : in    std_logic;
    P30CO   : out   std_logic;
    P30CTI  : in    std_logic;
    P30CTO  : out   std_logic;
    P30EI1  : in    std_logic;
    P30EI2  : in    std_logic;
    P30EI3  : in    std_logic;
    P30EI4  : in    std_logic;
    P30EI5  : in    std_logic;
    P30EI6  : in    std_logic;
    P30EI7  : in    std_logic;
    P30EI8  : in    std_logic;
    P30EL   : in    std_logic;
    P30ER   : in    std_logic;
    P30EO   : out   std_logic;
    P30RI   : in    std_logic;
    P30RL   : in    std_logic;
    P30RR   : in    std_logic;
    P30RO1  : out   std_logic;
    P30RO2  : out   std_logic;
    P30RO3  : out   std_logic;
    P30RO4  : out   std_logic;
    P30RO5  : out   std_logic;
    P30RO6  : out   std_logic;
    P30RO7  : out   std_logic;
    P30RO8  : out   std_logic;

    P31CI1  : in    std_logic;
    P31CL   : in    std_logic;
    P31CR   : in    std_logic;
    P31CO   : out   std_logic;
    P31CTI  : in    std_logic;
    P31CTO  : out   std_logic;
    P31EI1  : in    std_logic;
    P31EI2  : in    std_logic;
    P31EI3  : in    std_logic;
    P31EI4  : in    std_logic;
    P31EI5  : in    std_logic;
    P31EI6  : in    std_logic;
    P31EI7  : in    std_logic;
    P31EI8  : in    std_logic;
    P31EL   : in    std_logic;
    P31ER   : in    std_logic;
    P31EO   : out   std_logic;
    P31RI   : in    std_logic;
    P31RL   : in    std_logic;
    P31RR   : in    std_logic;
    P31RO1  : out   std_logic;
    P31RO2  : out   std_logic;
    P31RO3  : out   std_logic;
    P31RO4  : out   std_logic;
    P31RO5  : out   std_logic;
    P31RO6  : out   std_logic;
    P31RO7  : out   std_logic;
    P31RO8  : out   std_logic;

    P32CI1  : in    std_logic;
    P32CL   : in    std_logic;
    P32CR   : in    std_logic;
    P32CO   : out   std_logic;
    P32CTI  : in    std_logic;
    P32CTO  : out   std_logic;
    P32EI1  : in    std_logic;
    P32EI2  : in    std_logic;
    P32EI3  : in    std_logic;
    P32EI4  : in    std_logic;
    P32EI5  : in    std_logic;
    P32EI6  : in    std_logic;
    P32EI7  : in    std_logic;
    P32EI8  : in    std_logic;
    P32EL   : in    std_logic;
    P32ER   : in    std_logic;
    P32EO   : out   std_logic;
    P32RI   : in    std_logic;
    P32RL   : in    std_logic;
    P32RR   : in    std_logic;
    P32RO1  : out   std_logic;
    P32RO2  : out   std_logic;
    P32RO3  : out   std_logic;
    P32RO4  : out   std_logic;
    P32RO5  : out   std_logic;
    P32RO6  : out   std_logic;
    P32RO7  : out   std_logic;
    P32RO8  : out   std_logic;

    P33CI1  : in    std_logic;
    P33CL   : in    std_logic;
    P33CR   : in    std_logic;
    P33CO   : out   std_logic;
    P33CTI  : in    std_logic;
    P33CTO  : out   std_logic;
    P33EI1  : in    std_logic;
    P33EI2  : in    std_logic;
    P33EI3  : in    std_logic;
    P33EI4  : in    std_logic;
    P33EI5  : in    std_logic;
    P33EI6  : in    std_logic;
    P33EI7  : in    std_logic;
    P33EI8  : in    std_logic;
    P33EL   : in    std_logic;
    P33ER   : in    std_logic;
    P33EO   : out   std_logic;
    P33RI   : in    std_logic;
    P33RL   : in    std_logic;
    P33RR   : in    std_logic;
    P33RO1  : out   std_logic;
    P33RO2  : out   std_logic;
    P33RO3  : out   std_logic;
    P33RO4  : out   std_logic;
    P33RO5  : out   std_logic;
    P33RO6  : out   std_logic;
    P33RO7  : out   std_logic;
    P33RO8  : out   std_logic;

    P34CI1  : in    std_logic;
    P34CL   : in    std_logic;
    P34CR   : in    std_logic;
    P34CO   : out   std_logic;
    P34CTI  : in    std_logic;
    P34CTO  : out   std_logic;
    P34EI1  : in    std_logic;
    P34EI2  : in    std_logic;
    P34EI3  : in    std_logic;
    P34EI4  : in    std_logic;
    P34EI5  : in    std_logic;
    P34EI6  : in    std_logic;
    P34EI7  : in    std_logic;
    P34EI8  : in    std_logic;
    P34EL   : in    std_logic;
    P34ER   : in    std_logic;
    P34EO   : out   std_logic;
    P34RI   : in    std_logic;
    P34RL   : in    std_logic;
    P34RR   : in    std_logic;
    P34RO1  : out   std_logic;
    P34RO2  : out   std_logic;
    P34RO3  : out   std_logic;
    P34RO4  : out   std_logic;
    P34RO5  : out   std_logic;
    P34RO6  : out   std_logic;
    P34RO7  : out   std_logic;
    P34RO8  : out   std_logic
);
end NX_IOM_U;

-- =================================================================================================
--   NX_IOM_CONTROL_U definition                                                        2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_IOM_CONTROL_U is
generic (
    mode_side1        : integer := 0;
    div1         : bit_vector(2 downto 0) := "000";
    mode_side2        : integer := 0;
    div2         : bit_vector(2 downto 0) := "000";
    mode_side3        : integer := 0;
    div3         : bit_vector(2 downto 0) := "000";

    div_swrx1    : bit_vector(2 downto 0) := "000";
    div_swrx2    : bit_vector(2 downto 0) := "000";

    sel_ld_fck1  : bit_vector(1 downto 0) := "00";
    sel_ld_fck2  : bit_vector(1 downto 0) := "00";
    sel_ld_fck3  : bit_vector(1 downto 0) := "00";
    sel_sw_fck1  : bit_vector(1 downto 0) := "00";
    sel_sw_fck2  : bit_vector(1 downto 0) := "00";

    sel_dc_clk   : bit_vector(1 downto 0) := "00";

    inv_ld_sck1  : bit := '0';
    inv_ld_sck2  : bit := '0';
    inv_ld_sck3  : bit := '0';

    link_ld_12   : bit := '0';
    link_ld_23   : bit := '0';

    sel_clk_out1 : bit := '0';
    sel_clk_out2 : bit := '0';

    use_dc       : bit := '0';
    cal_delay1   : string := "";
    cal_delay2   : string := "";

    location     : string := ""
);
port(
    ALCK1   : in    std_logic;
    ALCK2   : in    std_logic;
    ALCK3   : in    std_logic;
    LDSCK1  : in    std_logic;
    LDSCK2  : in    std_logic;
    LDSCK3  : in    std_logic;
--  LDFCK1  : in    std_logic;	-- CONFIG
--  LDFCK2  : in    std_logic;	-- CONFIG
--  LDFCK3  : in    std_logic;	-- CONFIG
--  SWTX1CK : in    std_logic;	-- CONFIG
--  SWTX2CK : in    std_logic;	-- CONFIG
    SWRX1CK : in    std_logic;
    SWRX2CK : in    std_logic;
    FCK1    : in    std_logic;
    FCK2    : in    std_logic;
    FDCK    : in    std_logic;
    CCK     : in    std_logic;

    DQ1CI1  : in    std_logic;
    DQ1CI2  : in    std_logic;
    DQ1CI3  : in    std_logic;
    DQ1CI4  : in    std_logic;
    DQ1CI5  : in    std_logic;
    DQ1CI6  : in    std_logic;
    DQ1CI7  : in    std_logic;
    DQ1CI8  : in    std_logic;
    DQ2CI1  : in    std_logic;
    DQ2CI2  : in    std_logic;
    DQ2CI3  : in    std_logic;
    DQ2CI4  : in    std_logic;
    DQ2CI5  : in    std_logic;
    DQ2CI6  : in    std_logic;
    DQ2CI7  : in    std_logic;
    DQ2CI8  : in    std_logic;
    DQ3CI1  : in    std_logic;
    DQ3CI2  : in    std_logic;
    DQ3CI3  : in    std_logic;
    DQ3CI4  : in    std_logic;
    DQ3CI5  : in    std_logic;
    DQ3CI6  : in    std_logic;
    DQ3CI7  : in    std_logic;
    DQ3CI8  : in    std_logic;
    DQS1CI1 : in    std_logic;
    DQS1CI2 : in    std_logic;
    DQS1CI3 : in    std_logic;
    DQS1CI4 : in    std_logic;
    DQS1CI5 : in    std_logic;
    DQS1CI6 : in    std_logic;
    DQS1CI7 : in    std_logic;
    DQS1CI8 : in    std_logic;
    DQS2CI1 : in    std_logic;
    DQS2CI2 : in    std_logic;
    DQS2CI3 : in    std_logic;
    DQS2CI4 : in    std_logic;
    DQS2CI5 : in    std_logic;
    DQS2CI6 : in    std_logic;
    DQS2CI7 : in    std_logic;
    DQS2CI8 : in    std_logic;
    DQS3CI1 : in    std_logic;
    DQS3CI2 : in    std_logic;
    DQS3CI3 : in    std_logic;
    DQS3CI4 : in    std_logic;
    DQS3CI5 : in    std_logic;
    DQS3CI6 : in    std_logic;
    DQS3CI7 : in    std_logic;
    DQS3CI8 : in    std_logic;

    LD1RN   : in    std_logic;
    LD2RN   : in    std_logic;
    LD3RN   : in    std_logic;

    FA1     : in    std_logic;
    FA2     : in    std_logic;
    FA3     : in    std_logic;
    FA4     : in    std_logic;
    FA5     : in    std_logic;
    FA6     : in    std_logic;
    FZ      : in    std_logic;

    DCRN    : in    std_logic;
    LE      : in    std_logic;
    SE      : in    std_logic;

    DRI1     : in    std_logic;
    DRI2     : in    std_logic;
    DRI3     : in    std_logic;
    DRI4     : in    std_logic;
    DRI5     : in    std_logic;
    DRI6     : in    std_logic;
    DRA1     : in    std_logic;
    DRA2     : in    std_logic;
    DRA3     : in    std_logic;
    DRA4     : in    std_logic;

    DRO1CSN   : in    std_logic;
    DRO2CSN   : in    std_logic;
    DRO3CSN   : in    std_logic;
    DRI1CSN   : in    std_logic;
    DRI2CSN   : in    std_logic;
    DRI3CSN   : in    std_logic;
    DRDPA1CSN : in    std_logic;
    DRDPA2CSN : in    std_logic;
    DRDPA3CSN : in    std_logic;
    DRCCSN    : in    std_logic;
    DRWDS     : in    std_logic;
    DRWEN     : in    std_logic;
    DRE       : in    std_logic;

    CA1P1   : in    std_logic;
    CA1P2   : in    std_logic;
    CA1P3   : in    std_logic;
    CA1P4   : in    std_logic;
    CA2P1   : in    std_logic;
    CA2P2   : in    std_logic;
    CA2P3   : in    std_logic;
    CA2P4   : in    std_logic;
    CA1N1   : in    std_logic;
    CA1N2   : in    std_logic;
    CA1N3   : in    std_logic;
    CA1N4   : in    std_logic;
    CA2N1   : in    std_logic;
    CA2N2   : in    std_logic;
    CA2N3   : in    std_logic;
    CA2N4   : in    std_logic;
    CA1T1   : in    std_logic;
    CA1T2   : in    std_logic;
    CA1T3   : in    std_logic;
    CA1T4   : in    std_logic;
    CA2T1   : in    std_logic;
    CA2T2   : in    std_logic;
    CA2T3   : in    std_logic;
    CA2T4   : in    std_logic;
    CA1D1   : in    std_logic;
    CA1D2   : in    std_logic;
    CA1D3   : in    std_logic;
    CA1D4   : in    std_logic;
    CA1D5   : in    std_logic;
    CA1D6   : in    std_logic;
    CA2D1   : in    std_logic;
    CA2D2   : in    std_logic;
    CA2D3   : in    std_logic;
    CA2D4   : in    std_logic;
    CA2D5   : in    std_logic;
    CA2D6   : in    std_logic;

    CKO1    : out   std_logic;
    CKO2    : out   std_logic;

    FLD     : out   std_logic;
    FLG     : out   std_logic;
    AL1D    : out   std_logic;
    AL2D    : out   std_logic;
    AL3D    : out   std_logic;
    AL1T    : out   std_logic;
    AL2T    : out   std_logic;
    AL3T    : out   std_logic;
    DCL     : out   std_logic;
    DRO1    : out   std_logic;
    DRO2    : out   std_logic;
    DRO3    : out   std_logic;
    DRO4    : out   std_logic;
    DRO5    : out   std_logic;
    DRO6    : out   std_logic;

    LINK1  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK2  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK3  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK4  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK5  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK6  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK7  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK8  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK9  : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK10 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK11 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK12 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK13 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK14 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK15 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK16 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK17 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK18 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK19 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK20 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK21 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK22 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK23 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK24 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK25 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK26 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK27 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK28 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK29 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK30 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK31 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK32 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK33 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
    LINK34 : inout std_logic_vector(IOM_LINK_SIZE - 1 downto 0)
);
end NX_IOM_CONTROL_U;
-- =================================================================================================
--   NX_PLL_L definition                                                                2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

library NX;
use NX.nxPackage.all;

entity NX_PLL_L is
generic (
    location	      : string := "";
                      
    ref_intdiv        : integer   range 0 to 31 := 0;  -- 0 to 31  (%1 to %32)
    ref_osc_on        : bit := '0';                    -- 0: disabled - 1: enabled
                      
    cfg_use_pll       : std_logic:='1';                -- use or bypass PLL
                      
    ext_fbk_on        : bit := '0';                    -- 0: disabled - 1: enabled
                      
    fbk_intdiv        : integer   range 0 to 31 := 2;  -- 0 to 31  (%4 to %66 by step 2)
                      
    fbk_delay_on      : bit := '0';                    -- 0: no delay - 1: delay
    fbk_delay         : integer   range 0 to 63 := 0;  -- 0 to 63

    wfg_sync_pll_lock : bit := '0';                    -- 0: disabled - 1: enabled
    wfg_sync_cal_lock : bit := '0';                    -- 0: disabled - 1: enabled

    clk_outdivp1      : integer   range 0 to 7 := 0;   -- 0 to 7  P1 (2^n    : %1 to %128)
    clk_outdivp2      : integer   range 0 to 7 := 0;   -- 0 to 7  P2 (2^(n+1): %2 to %256)
    clk_outdivo1      : integer   range 0 to 7 := 0;   -- 0 to 7  O1 ((2n)+3 : %3 to  %17)
    clk_outdivp3o2    : integer   range 0 to 7 := 0    -- 0 to 7  P3 (2^(n+2): %4 to %512)
                                                       --         O2 ((2n)+5 : %5 to  %19)
);
port (
    REF               : in  std_logic;
    FBK               : in  std_logic;

    R                 : in  std_logic := '0';

    VCO               : out std_logic; -- CLK_PLL
    LDFO              : out std_logic; -- LDF_DIV
    REFO              : out std_logic; -- REF_DIV

    DIVO1             : out std_logic; -- (2n)+3
    DIVO2             : out std_logic; -- (2n)+5

    DIVP1             : out std_logic; -- 2^n
    DIVP2             : out std_logic; -- 2^(n+1)
    DIVP3             : out std_logic; -- 2^(n+2)
    OSC               : out std_logic; -- 100MHz

    PLL_LOCKED        : out std_logic;
    CAL_LOCKED        : out std_logic
);
end NX_PLL_L;

-- =================================================================================================
--   NX_WFG_L definition                                                                2018/11/30
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

library NX;
use NX.nxPackage.all;

entity NX_WFG_L is
generic (
    location    : string := "";
    wfg_edge    : bit := '0';                              -- 0: no invert / Rising
                                                           -- 1:    invert / Falling

    mode        : bit := '0';                              -- 0: no pattern - 1: pattern
    pattern_end : integer   range 0 to 15 := 1;            -- 0: to 15 (1 step to 16 steps)
    pattern     : bit_vector(0 to 15) := (others => '0');  -- pattern p0 ... p15

    delay_on    : bit := '0';                              -- 0: no delay - 1: delay
    delay       : integer   range 0 to 63 := 0             -- 0 to 63 (1 unit to 64 unit)
);
port (
    R   : in  std_logic := '0';
    SI  : in  std_logic;
    ZI  : in  std_logic;
    RDY : in  std_logic := '1';
    SO  : out std_logic;
    ZO  : out std_logic
);
end NX_WFG_L;

-- =================================================================================================
--   NX_PLL definition                                                                  2017/09/19
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

library NX;
use NX.nxPackage.all;

entity NX_PLL is
generic (
    location     : string := "";

    vco_range    : integer   range 0 to 2 := 0;   -- 0 to 3
    ref_div_on   : bit := '0';                    -- bypass :: %2
    fbk_div_on   : bit := '0';                    -- bypass :: %2
    ext_fbk_on   : bit := '0';                    -- 0: disabled - 1: enabled

    fbk_intdiv   : integer   range 1 to 31 := 2;  -- 0 to 31  (%1 to %32)

    fbk_delay_on : bit := '0';                    -- 0: no delay - 1: delay
    fbk_delay    : integer   range 0 to 63 := 0;  -- 0 to 63

    clk_outdiv1  : integer   range 0 to 7 := 0;   -- 0 to 7   (%1 to %2^7)
    clk_outdiv2  : integer   range 0 to 7 := 0;   -- 0 to 7   (%1 to %2^7)
    clk_outdiv3  : integer   range 0 to 7 := 0    -- 0 to 7   (%1 to %2^7)
);
port (
    REF : in  std_logic;
    FBK : in  std_logic;

    VCO : out std_logic;

    D1  : out std_logic;
    D2  : out std_logic;
    D3  : out std_logic;
    OSC : out std_logic;

    RDY : out std_logic
);
end NX_PLL;

-- =================================================================================================
--   NX_WFG definition                                                                  2017/09/19
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

library NX;
use NX.nxPackage.all;

entity NX_WFG is
generic (
    location    : string := "";

    wfg_edge    : bit := '0';                              -- 0: no invert / Rising
    mode        : bit := '0';                              -- 0: no pattern - 1: pattern

    pattern_end : integer   range 0 to 15 := 1;            -- 0: to 15 (1 step to 16 steps)
    pattern     : bit_vector(0 to 15) := (others => '0');  -- pattern p0 ... p15

    delay_on    : bit := '0';                              -- 0: no delay - 1: delay
    delay       : integer   range 0 to 63 := 0             -- 0 to 63 (1 unit to 64 unit)
);
port (
    SI  : in  std_logic;
    ZI  : in  std_logic;
    RDY : in  std_logic := '1';
    SO  : out std_logic;
    ZO  : out std_logic
);
end NX_WFG;

---------------------------------------------
--
-- NX_PLL_U.vhd
--
-- Creator : BEAU Sylvain
--
-- Editor : VSCode
--
-- 01/09/2020
---------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_PLL_U is
    generic (
        location     : string                 := "";               
        use_pll      : bit                    := '0';             -- Use the PLL
        pll_odf      : bit_vector(1 downto 0) := (others => '0'); -- Output division Factor
        pll_cpump    : bit_vector(3 downto 0) := (others => '0'); -- Set the charge pump factor
        pll_lpf_res  : bit_vector(3 downto 0) := (others => '0'); -- Set the resistances of the loop filter
        pll_lpf_cap  : bit_vector(3 downto 0) := (others => '0'); -- Set the capacitors of the loop filter
        pll_lock     : bit_vector(3 downto 0) := (others => '0'); -- Configuration of the frequency lock
        fbk_intdiv   : bit_vector(6 downto 0) := (others => '0'); -- Loop division Factor
        ref_intdiv   : bit_vector(4 downto 0) := (others => '0'); -- Reference Clock division Factor
        ref_osc_on   : bit                    := '0';             -- Reference Clock selection
        ext_fbk_on   : bit                    := '0';             -- Feedback Clock selection
        fbk_delay_on : bit                    := '0';             -- Add delay on the feedback clock
        fbk_delay    : bit_vector(5 downto 0) := (others => '0'); -- Delay on the feedback clock
        clk_outdiv1  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+3)
        clk_outdiv2  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+5)
        clk_outdiv3  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+7)
        clk_outdiv4  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (N+9)
        clk_outdivd1 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd2 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd3 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd4 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd5 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        use_cal      : bit                    := '0';             -- Use internal calibration
        clk_cal_sel  : bit_vector(1 downto 0) := "01";            -- Internal calibration clock selector
        cal_div      : bit_vector(3 downto 0) := "0111";          -- Division factor on Internal calibration clock
        cal_delay    : bit_vector(5 downto 0) := "011011"         -- Delay on internal calibration clock
    );
    port (
        R              : in std_logic;  -- Reset
        REF            : in std_logic;  -- PLL's reference clock
        FBK            : in std_logic;  -- PLL's feedback clock
        -- Clock
        OSC            : out std_logic; -- Oscillator's clock
        VCO            : out std_logic; -- PLL's output
        LDFO           : out std_logic; -- LDF_DIV
        REFO           : out std_logic; -- REF_DIV
        CLK_DIV1       : out std_logic; -- 1/(N+3)
        CLK_DIV2       : out std_logic; -- 1/(N+5)
        CLK_DIV3       : out std_logic; -- 1/(N+7)
        CLK_DIV4       : out std_logic; -- 1/(N+9)
        CLK_DIVD1     : out std_logic; -- 1/(N+2)
        CLK_DIVD2     : out std_logic; -- 1/(N+2)
        CLK_DIVD3     : out std_logic; -- 1/(N+2)
        CLK_DIVD4     : out std_logic; -- 1/(N+2)
        CLK_DIVD5     : out std_logic; -- 1/(N+2)
        -- Lock engine
        PLL_LOCKED     : out std_logic;
        PLL_LOCKEDA    : out std_logic;
        -- Calbration
        ARST_CAL       : in std_logic;  -- calibration's reset
        CLK_CAL        : in std_logic;  -- Calibration's clock
        CLK_CAL_DIV    : out std_logic; -- Output of calibration clock's divider
        CAL_LOCKED     : out std_logic;
        EXT_CAL_LOCKED : in std_logic;
        CAL1           : out std_logic;
        CAL2           : out std_logic;
        CAL3           : out std_logic;
        CAL4           : out std_logic;
        CAL5           : out std_logic;
        EXT_CAL1       : in std_logic;
        EXT_CAL2       : in std_logic;
        EXT_CAL3       : in std_logic;
        EXT_CAL4       : in std_logic;
        EXT_CAL5       : in std_logic
    );
end NX_PLL_U;
---------------------------------------------
--
-- NX_PLL_U_WRAPPER.vhd
--
-- Creator : BEAU Sylvain
--
-- Editor : VSCode
--
-- 01/09/2020
---------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity NX_PLL_U_WRAP is
    generic (
        location     : string                 := ""; 
        use_pll      : bit                    := '0';             -- Use the PLL
        pll_odf      : bit_vector(1 downto 0) := (others => '0'); -- Output division Factor
        pll_cpump    : bit_vector(3 downto 0) := (others => '0'); -- Set the charge pump factor
        pll_lpf_res  : bit_vector(3 downto 0) := (others => '0'); -- Set the resistances of the loop filter
        pll_lpf_cap  : bit_vector(3 downto 0) := (others => '0'); -- Set the capacitors of the loop filter
        pll_lock     : bit_vector(3 downto 0) := (others => '0'); -- Configuration of the frequency lock
        fbk_intdiv   : bit_vector(6 downto 0) := (others => '0'); -- Loop division Factor
        ref_intdiv   : bit_vector(4 downto 0) := (others => '0'); -- Reference Clock division Factor
        ref_osc_on   : bit                    := '0';             -- Reference Clock selection
        ext_fbk_on   : bit                    := '0';             -- Feedback Clock selection
        fbk_delay_on : bit                    := '0';             -- Add delay on the feedback clock
        fbk_delay    : bit_vector(5 downto 0) := (others => '0'); -- Delay on the feedback clock
        clk_outdiv1  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+3)
        clk_outdiv2  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+5)
        clk_outdiv3  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+7)
        clk_outdiv4  : bit_vector(2 downto 0) := (others => '0'); -- PLL division Factor (2*N+9)
        clk_outdivd1 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd2 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd3 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd4 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        clk_outdivd5 : bit_vector(3 downto 0) := (others => '0'); -- PLL division Factor (N+2)
        use_cal      : bit                    := '0';             -- Use internal calibration
        clk_cal_sel  : bit_vector(1 downto 0) := "01";            -- Internal calibration clock selector
        cal_div      : bit_vector(3 downto 0) := "0111";          -- Division factor on Internal calibration clock
        cal_delay    : bit_vector(5 downto 0) := "011011"         -- Delay on internal calibration clock
    );
    port (
        R              : in std_logic;  -- Reset
        REF            : in std_logic;  -- PLL's reference clock
        FBK            : in std_logic;  -- PLL's feedback clock
        -- Clock
        OSC            : out std_logic; -- Oscillator's clock
        VCO            : out std_logic; -- PLL's output
        LDFO           : out std_logic; -- LDF_DIV
        REFO           : out std_logic; -- REF_DIV
        CLK_DIV        : out std_logic_vector(3 downto 0); -- 0 : 1/(N+3); 1 : 1/(N+5); 2 : 1/(N+7); 3 : 1/(N+9)
        CLK_DIVD       : out std_logic_vector(4 downto 0); -- 1/(N+2)
        -- Lock engine
        PLL_LOCKED     : out std_logic;
        PLL_LOCKEDA    : out std_logic;
        -- Calibration
        ARST_CAL       : in std_logic;  -- calibration's reset
        CLK_CAL        : in std_logic;  -- calibration's clock
        CLK_CAL_DIV    : out std_logic;
        CAL_LOCKED     : out std_logic;
        EXT_CAL_LOCKED : in std_logic;
        CAL            : out std_logic_vector(4 downto 0);
        EXT_CAL        : in std_logic_vector(4 downto 0)
    );
end NX_PLL_U_WRAP;

architecture NX_RTL of NX_PLL_U_WRAP is

    component NX_PLL_U
        generic (
	     location     : string                := "";--  
            use_pll      : bit                    := '0';--
            pll_odf      : bit_vector(1 downto 0) := (others => '0');--
            pll_cpump    : bit_vector(3 downto 0) := (others => '0');--
            pll_lpf_res  : bit_vector(3 downto 0) := (others => '0');--
            pll_lpf_cap  : bit_vector(3 downto 0) := (others => '0');--
            pll_lock     : bit_vector(3 downto 0) := (others => '0');
            fbk_intdiv   : bit_vector(6 downto 0) := (others => '0');--
            ref_intdiv   : bit_vector(4 downto 0) := (others => '0');--
            ref_osc_on   : bit                    := '0';--
            ext_fbk_on   : bit                    := '0';--
            fbk_delay_on : bit                    := '0';--
            fbk_delay    : bit_vector(5 downto 0) := (others => '0');--
            clk_outdiv1  : bit_vector(2 downto 0) := (others => '0');--
            clk_outdiv2  : bit_vector(2 downto 0) := (others => '0');--
            clk_outdiv3  : bit_vector(2 downto 0) := (others => '0');--
            clk_outdiv4  : bit_vector(2 downto 0) := (others => '0');--
            clk_outdivd1 : bit_vector(3 downto 0) := (others => '0');--
            clk_outdivd2 : bit_vector(3 downto 0) := (others => '0');--
            clk_outdivd3 : bit_vector(3 downto 0) := (others => '0');--
            clk_outdivd4 : bit_vector(3 downto 0) := (others => '0');--
            clk_outdivd5 : bit_vector(3 downto 0) := (others => '0');--
            use_cal      : bit                    := '0';
            clk_cal_sel  : bit_vector(1 downto 0) := "01";
            cal_div      : bit_vector(3 downto 0) := "0111";
            cal_delay    : bit_vector(5 downto 0) := "011011"
        );
        port (
            OSC            : out std_logic;--
            REF            : in std_logic;--
            FBK            : in std_logic;--
            R              : in std_logic;--
            CLK_CAL        : in std_logic;
            VCO            : out std_logic;--
            LDFO           : out std_logic;--
            REFO           : out std_logic;--
            CLK_DIV1       : out std_logic;
            CLK_DIV2       : out std_logic;
            CLK_DIV3       : out std_logic;
            CLK_DIV4       : out std_logic;
            CLK_DIVD1      : out std_logic;--
            CLK_DIVD2      : out std_logic;--
            CLK_DIVD3      : out std_logic;--
            CLK_DIVD4      : out std_logic;--
            CLK_DIVD5      : out std_logic;--
            PLL_LOCKED     : out std_logic;--
            PLL_LOCKEDA    : out std_logic;
            ARST_CAL       : in std_logic;--
            CLK_CAL_DIV    : out std_logic;--
            CAL_LOCKED     : out std_logic;--
            EXT_CAL_LOCKED : in std_logic;--
            CAL1           : out std_logic;--
            CAL2           : out std_logic;--
            CAL3           : out std_logic;--
            CAL4           : out std_logic;--
            CAL5           : out std_logic;--
            EXT_CAL1       : in std_logic;
            EXT_CAL2       : in std_logic;
            EXT_CAL3       : in std_logic;
            EXT_CAL4       : in std_logic;
            EXT_CAL5       : in std_logic --
        );
    end component;

begin

    pll : NX_PLL_U
    generic map (
        location     => location,     -- string             := "";
        use_pll      => use_pll,      -- bit                := '0';--
        pll_odf      => pll_odf,      -- bit_vector(0 to 1) := (others => '0');--
        pll_cpump    => pll_cpump,    -- bit_vector(0 to 3) := (others => '0');--
        pll_lpf_res  => pll_lpf_res,  -- bit_vector(0 to 3) := (others => '0');--
        pll_lpf_cap  => pll_lpf_cap,  -- bit_vector(0 to 3) := (others => '0');--
        pll_lock     => pll_lock,     -- bit_vector(0 to 3) := (others => '0');
        fbk_intdiv   => fbk_intdiv,   -- bit_vector(0 to 6) := (others => '0');--
        ref_intdiv   => ref_intdiv,   -- bit_vector(0 to 4) := (others => '0');--
        ref_osc_on   => ref_osc_on,   -- bit                := '0';--
        ext_fbk_on   => ext_fbk_on,   -- bit                := '0';--
        fbk_delay_on => fbk_delay_on, -- bit                := '0';--
        fbk_delay    => fbk_delay,    -- bit_vector(0 to 5) := (others => '0');--
        clk_outdiv1  => clk_outdiv1,  -- bit_vector(0 to 2) := (others => '0');--
        clk_outdiv2  => clk_outdiv2,  -- bit_vector(0 to 2) := (others => '0');--
        clk_outdiv3  => clk_outdiv3,  -- bit_vector(0 to 2) := (others => '0');--
        clk_outdiv4  => clk_outdiv4,  -- bit_vector(0 to 2) := (others => '0');--
        clk_outdivd1 => clk_outdivd1, -- bit_vector(0 to 3) := (others => '0');--
        clk_outdivd2 => clk_outdivd2, -- bit_vector(0 to 3) := (others => '0');--
        clk_outdivd3 => clk_outdivd3, -- bit_vector(0 to 3) := (others => '0');--
        clk_outdivd4 => clk_outdivd4, -- bit_vector(0 to 3) := (others => '0');--
        clk_outdivd5 => clk_outdivd5, -- bit_vector(0 to 3) := (others => '0');--
        use_cal      => use_cal,      -- bit                := '0';
        clk_cal_sel  => clk_cal_sel,  -- bit_vector(0 to 1) := "01";
        cal_div      => cal_div,      -- bit_vector(0 to 3) := "0111";
        cal_delay    => cal_delay     -- bit_vector(0 to 5) := "011011"
    )
    port map (
        OSC            => OSC, -- out std_logic;--
        REF            => REF, -- in std_logic;--
        FBK            => FBK, -- in std_logic;--
        R              => R, -- in std_logic;--
        CLK_CAL        => CLK_CAL, -- in std_logic;
        VCO            => VCO, -- out std_logic;--
        LDFO           => LDFO, -- out std_logic;--
        REFO           => REFO, -- out std_logic;--
        CLK_DIV1       => CLK_DIV(0), -- out std_logic;
        CLK_DIV2       => CLK_DIV(1), -- out std_logic;
        CLK_DIV3       => CLK_DIV(2), -- out std_logic;
        CLK_DIV4       => CLK_DIV(3), -- out std_logic;
        CLK_DIVD1      => CLK_DIVD(0), -- out std_logic;--
        CLK_DIVD2      => CLK_DIVD(1), -- out std_logic;--
        CLK_DIVD3      => CLK_DIVD(2), -- out std_logic;--
        CLK_DIVD4      => CLK_DIVD(3), -- out std_logic;--
        CLK_DIVD5      => CLK_DIVD(4), -- out std_logic;--
        PLL_LOCKED     => PLL_LOCKED, -- out std_logic;--
        PLL_LOCKEDA    => PLL_LOCKEDA, -- out std_logic;
        ARST_CAL       => ARST_CAL, -- in std_logic;--
        CLK_CAL_DIV    => CLK_CAL_DIV, -- out std_logic;--
        CAL_LOCKED     => CAL_LOCKED, -- out std_logic;--
        EXT_CAL_LOCKED => EXT_CAL_LOCKED, -- in std_logic;--
        CAL1           => CAL(0), -- out std_logic;--
        CAL2           => CAL(1), -- out std_logic;--
        CAL3           => CAL(2), -- out std_logic;--
        CAL4           => CAL(3), -- out std_logic;--
        CAL5           => CAL(4), -- out std_logic;--
        EXT_CAL1       => EXT_CAL(0), -- in std_logic;
        EXT_CAL2       => EXT_CAL(1), -- in std_logic;
        EXT_CAL3       => EXT_CAL(2), -- in std_logic;
        EXT_CAL4       => EXT_CAL(3), -- in std_logic;
        EXT_CAL5       => EXT_CAL(4)  -- in std_logic;--
    );

end NX_RTL;
---------------------------------------------
--
-- NX_WFG_U.vhd
--
-- Creator : BEAU Sylvain
--
-- Editor : VSCode
--
-- 01/09/2020
---------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library NX;
use NX.nxPackage.all;

entity NX_WFG_U is
    generic (
        location             : string := "";
        wfg_edge             : bit                   := '0'; -- 0: no invert / Rising
        reset_on_pll_lock_n  : bit                   := '0';
        reset_on_pll_locka_n : bit                   := '0';
        reset_on_cal_lock_n  : bit                   := '0';

        mode                 : integer range 0 to 2 := 0;                                   -- 0: no pattern - 1: pattern - 2: diviseur
        pattern              : bit_vector(0 to 15)   := b"0000000000000000"; -- pattern p0 ... p15
        pattern_end          : integer range 0 to 15 := 0;                   -- max pattern length. Set to 0 to use divider/bypass instead of pattern
        div_ratio            : integer range 0 to 2047 := 0;                   -- divisor ratio
        delay_on             : bit                   := '0';                 -- 0: no delay - 1: delay
        delay                : integer range 0 to 63 := 0                    -- 0 to 63 (1 unit to 32 unit)
    );
    port (
        R  : in std_logic;
        SI : in std_logic;
        ZI : in std_logic;
        SO : out std_logic;
        ZO : out std_logic
    );
end NX_WFG_U;
-- =================================================================================================
--   NX_R5_L definition                                                                 2019/04/09
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_R5_L is
port (
    -- Inputs
    A_CKEM_I      : in  std_logic; --  aclkenm0      1
    A_CKEP_I      : in  std_logic; --  aclkenp0      1
    A_CKES_I      : in  std_logic; --  aclkens0      1

    AR_A_I32      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I31      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I30      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I29      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I28      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I27      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I26      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I25      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I24      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I23      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I22      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I21      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I20      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I19      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I18      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I17      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I16      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I15      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I14      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I13      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I12      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I11      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I10      : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I9       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I8       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I7       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I6       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I5       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I4       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I3       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I2       : in  std_logic; --  araddrs0      32  [0:31]
    AR_A_I1       : in  std_logic; --  araddrs0      32  [0:31]

    AR_BU_I2      : in  std_logic; --  arbursts0     2   [0:1]
    AR_BU_I1      : in  std_logic; --  arbursts0     2   [0:1]

    AR_CH_I4      : in  std_logic; --  arcaches0     4   [0:3]
    AR_CH_I3      : in  std_logic; --  arcaches0     4   [0:3]
    AR_CH_I2      : in  std_logic; --  arcaches0     4   [0:3]
    AR_CH_I1      : in  std_logic; --  arcaches0     4   [0:3]

    AR_IDS_I8     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I7     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I6     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I5     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I4     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I3     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I2     : in  std_logic; --  arids0        8   [0:7]
    AR_IDS_I1     : in  std_logic; --  arids0        8   [0:7]

    AR_LE_I4      : in  std_logic; --  arlens0       4   [0:3]
    AR_LE_I3      : in  std_logic; --  arlens0       4   [0:3]
    AR_LE_I2      : in  std_logic; --  arlens0       4   [0:3]
    AR_LE_I1      : in  std_logic; --  arlens0       4   [0:3]

    AR_LK_I2      : in  std_logic; --  arlocks0      2   [0:1]
    AR_LK_I1      : in  std_logic; --  arlocks0      2   [0:1]

    AR_PR_I3      : in  std_logic; --  arprots0      3   [0:2]
    AR_PR_I2      : in  std_logic; --  arprots0      3   [0:2]
    AR_PR_I1      : in  std_logic; --  arprots0      3   [0:2]

    AR_RYM_I      : in  std_logic; --  arreadym0     1
    AR_RYP_I      : in  std_logic; --  arreadyp0     1

    AR_SZ_I3      : in  std_logic; --  arsizes0      3   [0:2]
    AR_SZ_I2      : in  std_logic; --  arsizes0      3   [0:2]
    AR_SZ_I1      : in  std_logic; --  arsizes0      3   [0:2]

    AR_VD_I       : in  std_logic; --  arvalids0     1
    AT_RS_I       : in  std_logic; --  atresetn      1

    AW_A_I32      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I31      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I30      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I29      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I28      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I27      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I26      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I25      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I24      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I23      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I22      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I21      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I20      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I19      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I18      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I17      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I16      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I15      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I14      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I13      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I12      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I11      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I10      : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I9       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I8       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I7       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I6       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I5       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I4       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I3       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I2       : in  std_logic; --  awaddrs0      32  [0:31]
    AW_A_I1       : in  std_logic; --  awaddrs0      32  [0:31]

    AW_BU_I2      : in  std_logic; --  awbursts0     2   [0:1]
    AW_BU_I1      : in  std_logic; --  awbursts0     2   [0:1]

    AW_CH_I4      : in  std_logic; --  awcaches0     4   [0:3]
    AW_CH_I3      : in  std_logic; --  awcaches0     4   [0:3]
    AW_CH_I2      : in  std_logic; --  awcaches0     4   [0:3]
    AW_CH_I1      : in  std_logic; --  awcaches0     4   [0:3]

    AW_IDS_I8     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I7     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I6     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I5     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I4     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I3     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I2     : in  std_logic; --  awids0        8   [0:7]
    AW_IDS_I1     : in  std_logic; --  awids0        8   [0:7]

    AW_LE_I4      : in  std_logic; --  awlens0       4   [0:3]
    AW_LE_I3      : in  std_logic; --  awlens0       4   [0:3]
    AW_LE_I2      : in  std_logic; --  awlens0       4   [0:3]
    AW_LE_I1      : in  std_logic; --  awlens0       4   [0:3]

    AW_LK_I2      : in  std_logic; --  awlocks0      2   [0:1]
    AW_LK_I1      : in  std_logic; --  awlocks0      2   [0:1]

    AW_PR_I3      : in  std_logic; --  awprots0      3   [0:2]
    AW_PR_I2      : in  std_logic; --  awprots0      3   [0:2]
    AW_PR_I1      : in  std_logic; --  awprots0      3   [0:2]

    AW_RYM_I      : in  std_logic; --  awreadym0     1
    AW_RYP_I      : in  std_logic; --  awreadyp0     1

    AW_SZ_I3      : in  std_logic; --  awsizes0      3   [0:2]
    AW_SZ_I2      : in  std_logic; --  awsizes0      3   [0:2]
    AW_SZ_I1      : in  std_logic; --  awsizes0      3   [0:2]

    AW_VD_I       : in  std_logic; --  awvalids0     1

    B_IDM_I4      : in  std_logic; --  bidm0         4   [0:3]
    B_IDM_I3      : in  std_logic; --  bidm0         4   [0:3]
    B_IDM_I2      : in  std_logic; --  bidm0         4   [0:3]
    B_IDM_I1      : in  std_logic; --  bidm0         4   [0:3]

    B_IDP_I4      : in  std_logic; --  bidp0         4   [0:3]
    B_IDP_I3      : in  std_logic; --  bidp0         4   [0:3]
    B_IDP_I2      : in  std_logic; --  bidp0         4   [0:3]
    B_IDP_I1      : in  std_logic; --  bidp0         4   [0:3]

    B_RDY_I       : in  std_logic; --  breadys0      1

    B_RSPM_I2     : in  std_logic; --  brespm0 2     [0:1]
    B_RSPM_I1     : in  std_logic; --  brespm0 2     [0:1]

    B_RSPP_I2     : in  std_logic; --  brespp0 2     [0:1]
    B_RSPP_I1     : in  std_logic; --  brespp0 2     [0:1]

    B_VDM_I       : in  std_logic; --  bvalidm0      1
    B_VDP_I       : in  std_logic; --  bvalidp0      1

--    CAL_I5        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I4        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I3        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I2        : in  std_logic; --  calibration   5   [0:4]
--    CAL_I1        : in  std_logic; --  calibration   5   [0:4]

    CDB_PW_I      : in  std_logic; --  cdbgpwrupack  1
    CDB_RS_I      : in  std_logic; --  cdbgrstack    1
    CFG_EE_I      : in  std_logic; --  cfgee         1
    CFG_IE_I      : in  std_logic; --  cfgie         1
    CFG_NM_I      : in  std_logic; --  cfgnmfi0      1
    CK_I          : in  std_logic; --  clk           1
--    CK_DR_I       : in  std_logic; --  clock_dr      1
    CS_PW_I       : in  std_logic; --  csyspwrupack  1
    DB_E_I        : in  std_logic; --  dbgen0        1
    DB_NCK_I      : in  std_logic; --  dbgnoclkstop  1

    DB_RA_I20     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I19     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I18     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I17     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I16     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I15     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I14     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I13     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I12     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I11     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I10     : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I9      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I8      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I7      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I6      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I5      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I4      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I3      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I2      : in  std_logic; --  dbgromaddr    20  [0:19]
    DB_RA_I1      : in  std_logic; --  dbgromaddr    20  [0:19]

    DB_RAV_I      : in  std_logic; --  dbgromaddrv   1

    DB_SA_I20     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I19     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I18     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I17     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I16     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I15     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I14     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I13     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I12     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I11     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I10     : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I9      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I8      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I7      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I6      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I5      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I4      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I3      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I2      : in  std_logic; --  dbgselfaddr0  20  [0:19]
    DB_SA_I1      : in  std_logic; --  dbgselfaddr0  20  [0:19]

    DB_SAV_I      : in  std_logic; --  dbgselfaddrv0 1
    DEV_E_I       : in  std_logic; --  deviceen      1

    DFTS_I8       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I7       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I6       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I5       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I4       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I3       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I2       : in  std_logic; --  dftsi         8   [0:7]
    DFTS_I1       : in  std_logic; --  dftsi         8   [0:7]

    E_DB_I        : in  std_logic; --  edbgrq0       1
    ERR_R_I       : in  std_logic; --  errenram0     1
    EVENT_I       : in  std_logic; --  eventi0       1

    GID_I4        : in  std_logic; --  groupid       4   [0:3]
    GID_I3        : in  std_logic; --  groupid       4   [0:3]
    GID_I2        : in  std_logic; --  groupid       4   [0:3]
    GID_I1        : in  std_logic; --  groupid       4   [0:3]

    INIT_P_I      : in  std_logic; --  initppx0      1
    INIT_R_I      : in  std_logic; --  initrama0     1
    LOC_R_I       : in  std_logic; --  loczrama0     1
--    LBK_E_I       : in  std_logic; --  loopback_en   1
--    LBK_MX_I      : in  std_logic; --  loopback_mux  1

--    MODE1_I3      : in  std_logic; --  mode1         3   [0:2]
--    MODE1_I2      : in  std_logic; --  mode1         3   [0:2]
--    MODE1_I1      : in  std_logic; --  mode1         3   [0:2]

--    MODE2_I3      : in  std_logic; --  mode2         3   [0:2]
--    MODE2_I2      : in  std_logic; --  mode2         3   [0:2]
--    MODE2_I1      : in  std_logic; --  mode2         3   [0:2]

--    MODE3_I3      : in  std_logic; --  mode3         3   [0:2]
--    MODE3_I2      : in  std_logic; --  mode3         3   [0:2]
--    MODE3_I1      : in  std_logic; --  mode3         3   [0:2]

    NCPUH_I       : in  std_logic; --  ncpuhalt0     1
    NET_RS_I      : in  std_logic; --  netmporeset   1
    N_FIQ_I       : in  std_logic; --  nfiq0         1
    N_IDE_I       : in  std_logic; --  niden0        1
    N_IRQ_I       : in  std_logic; --  nirq0         1
    N_PRS_I       : in  std_logic; --  npotrst       1
    N_RS_I        : in  std_logic; --  nreset0       1
    N_SPRS_I      : in  std_logic; --  nsysporeset   1
    N_TRS_I       : in  std_logic; --  ntrst         1

    P_A_I29       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I28       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I27       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I26       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I25       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I24       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I23       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I22       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I21       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I20       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I19       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I18       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I17       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I16       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I15       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I14       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I13       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I12       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I11       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I10       : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I9        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I8        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I7        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I6        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I5        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I4        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I3        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I2        : in  std_logic; --  paddrsys      29  [0:28]
    P_A_I1        : in  std_logic; --  paddrsys      29  [0:28]

    P_ECC_I       : in  std_logic; --  pareccenram0  1
    PLVL_I        : in  std_logic; --  paritylevel   1
    P_CK_E_I      : in  std_logic; --  pclkensys     1
    P_CK_I        : in  std_logic; --  pclksys       1
    P_E_I         : in  std_logic; --  penablesys    1

    PPV_BS_I20    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I19    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I18    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I17    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I16    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I15    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I14    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I13    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I12    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I11    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I10    : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I9     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I8     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I7     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I6     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I5     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I4     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I3     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I2     : in  std_logic; --  ppvbase0      20  [0:19]
    PPV_BS_I1     : in  std_logic; --  ppvbase0      20  [0:19]

    PPV_SZ_I5     : in  std_logic; --  ppvsize0      5   [0:4]
    PPV_SZ_I4     : in  std_logic; --  ppvsize0      5   [0:4]
    PPV_SZ_I3     : in  std_logic; --  ppvsize0      5   [0:4]
    PPV_SZ_I2     : in  std_logic; --  ppvsize0      5   [0:4]
    PPV_SZ_I1     : in  std_logic; --  ppvsize0      5   [0:4]

    PPX_BS_I20    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I19    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I18    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I17    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I16    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I15    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I14    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I13    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I12    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I11    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I10    : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I9     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I8     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I7     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I6     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I5     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I4     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I3     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I2     : in  std_logic; --  ppxbase0      20  [0:19]
    PPX_BS_I1     : in  std_logic; --  ppxbase0      20  [0:19]

    PPX_SZ_I5     : in  std_logic; --  ppxsize0      5   [0:4]
    PPX_SZ_I4     : in  std_logic; --  ppxsize0      5   [0:4]
    PPX_SZ_I3     : in  std_logic; --  ppxsize0      5   [0:4]
    PPX_SZ_I2     : in  std_logic; --  ppxsize0      5   [0:4]
    PPX_SZ_I1     : in  std_logic; --  ppxsize0      5   [0:4]

    P_RS_I        : in  std_logic; --  presetsysn    1
    P_SEL_I       : in  std_logic; --  pselsys       1

    PW_D_I32      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I31      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I30      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I29      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I28      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I27      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I26      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I25      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I24      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I23      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I22      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I21      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I20      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I19      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I18      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I17      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I16      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I15      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I14      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I13      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I12      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I11      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I10      : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I9       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I8       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I7       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I6       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I5       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I4       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I3       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I2       : in  std_logic; --  pwdatasys     32  [0:31]
    PW_D_I1       : in  std_logic; --  pwdatasys     32  [0:31]

    PW_I          : in  std_logic; --  pwritesys     1

    RAMCTL_I8     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I7     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I6     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I5     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I4     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I3     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I2     : in  std_logic; --  ramcontrol0   8   [0:7]
    RAMCTL_I1     : in  std_logic; --  ramcontrol0   8   [0:7]

    R_DM_I64      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I63      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I62      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I61      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I60      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I59      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I58      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I57      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I56      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I55      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I54      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I53      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I52      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I51      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I50      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I49      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I48      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I47      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I46      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I45      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I44      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I43      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I42      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I41      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I40      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I39      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I38      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I37      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I36      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I35      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I34      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I33      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I32      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I31      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I30      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I29      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I28      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I27      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I26      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I25      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I24      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I23      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I22      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I21      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I20      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I19      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I18      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I17      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I16      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I15      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I14      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I13      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I12      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I11      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I10      : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I9       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I8       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I7       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I6       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I5       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I4       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I3       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I2       : in  std_logic; --  rdatam0       64  [0:63]
    R_DM_I1       : in  std_logic; --  rdatam0       64  [0:63]

    R_DP_I32      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I31      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I30      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I29      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I28      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I27      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I26      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I25      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I24      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I23      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I22      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I21      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I20      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I19      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I18      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I17      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I16      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I15      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I14      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I13      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I12      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I11      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I10      : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I9       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I8       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I7       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I6       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I5       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I4       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I3       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I2       : in  std_logic; --  rdatap0       32  [0:31]
    R_DP_I1       : in  std_logic; --  rdatap0       32  [0:31]

--    RDY_I3        : in  std_logic; --  ready         3   [0:2]
--    RDY_I2        : in  std_logic; --  ready         3   [0:2]
--    RDY_I1        : in  std_logic; --  ready         3   [0:2]

    R_IDM_I4      : in  std_logic; --  ridm0         4   [0:3]
    R_IDM_I3      : in  std_logic; --  ridm0         4   [0:3]
    R_IDM_I2      : in  std_logic; --  ridm0         4   [0:3]
    R_IDM_I1      : in  std_logic; --  ridm0         4   [0:3]

    R_IDP_I4      : in  std_logic; --  ridp0         4   [0:3]
    R_IDP_I3      : in  std_logic; --  ridp0         4   [0:3]
    R_IDP_I2      : in  std_logic; --  ridp0         4   [0:3]
    R_IDP_I1      : in  std_logic; --  ridp0         4   [0:3]

    R_LSTM_I      : in  std_logic; --  rlastm0       1
    R_LSTP_I      : in  std_logic; --  rlastp0       1
    R_RDY_I       : in  std_logic; --  rreadys0      1

    R_RSPM_I2     : in  std_logic; --  rrespm0       2   [0:1]
    R_RSPM_I1     : in  std_logic; --  rrespm0       2   [0:1]

    R_RSPP_I2     : in  std_logic; --  rrespp0       2   [0:1]
    R_RSPP_I1     : in  std_logic; --  rrespp0       2   [0:1]

    RS_BYP_I      : in  std_logic; --  rstbypass     1
    R_VDM_I       : in  std_logic; --  rvalidm0      1
    R_VDP_I       : in  std_logic; --  rvalidp0      1
--    SCAN_E_I      : in  std_logic; --  scan_en       1
    SE_I          : in  std_logic; --  se            1
--    SHF_DR_I      : in  std_logic; --  shift_dr      1
--    SH_I          : in  std_logic; --  shin          1
    SW_CK_I       : in  std_logic; --  swclktck      1
    SW_DI_I       : in  std_logic; --  swditms       1
    T_DI_I        : in  std_logic; --  tdi           1
    TE_INI_I      : in  std_logic; --  teinit        1
--    TEST_E_I      : in  std_logic; --  test_en       1
--    UPD_DR_I      : in  std_logic; --  update_dr     1
    VINI_I        : in  std_logic; --  vinithi0      1

    W_D_I64       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I63       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I62       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I61       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I60       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I59       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I58       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I57       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I56       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I55       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I54       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I53       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I52       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I51       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I50       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I49       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I48       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I47       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I46       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I45       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I44       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I43       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I42       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I41       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I40       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I39       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I38       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I37       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I36       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I35       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I34       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I33       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I32       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I31       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I30       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I29       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I28       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I27       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I26       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I25       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I24       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I23       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I22       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I21       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I20       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I19       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I18       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I17       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I16       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I15       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I14       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I13       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I12       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I11       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I10       : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I9        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I8        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I7        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I6        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I5        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I4        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I3        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I2        : in  std_logic; --  wdatas0       64  [0:63]
    W_D_I1        : in  std_logic; --  wdatas0       64  [0:63]

    W_IDS_I8      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I7      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I6      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I5      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I4      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I3      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I2      : in  std_logic; --  wids0         8   [0:7]
    W_IDS_I1      : in  std_logic; --  wids0         8   [0:7]

    W_LST_I       : in  std_logic; --  wlasts0       1
    W_RYM_I       : in  std_logic; --  wreadym0      1
    W_RYP_I       : in  std_logic; --  wreadyp0      1

    W_SBS_I8      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I7      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I6      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I5      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I4      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I3      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I2      : in  std_logic; --  wstrbs0       8   [0:7]
    W_SBS_I1      : in  std_logic; --  wstrbs0       8   [0:7]

    W_VD_I        : in  std_logic; --  wvalids0      1

    -- Outputs
    AR_AM_O32     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O31     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O30     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O29     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O28     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O27     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O26     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O25     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O24     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O23     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O22     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O21     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O20     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O19     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O18     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O17     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O16     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O15     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O14     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O13     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O12     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O11     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O10     : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O9      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O8      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O7      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O6      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O5      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O4      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O3      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O2      : out std_logic; --  araddrm0            32  [0:31]
    AR_AM_O1      : out std_logic; --  araddrm0            32  [0:31]

    AR_AP_O32     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O31     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O30     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O29     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O28     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O27     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O26     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O25     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O24     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O23     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O22     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O21     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O20     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O19     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O18     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O17     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O16     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O15     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O14     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O13     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O12     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O11     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O10     : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O9      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O8      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O7      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O6      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O5      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O4      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O3      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O2      : out std_logic; --  araddrp0            32  [0:31]
    AR_AP_O1      : out std_logic; --  araddrp0            32  [0:31]

    AR_BUM_O2     : out std_logic; --  arburstm0           2   [0:1]
    AR_BUM_O1     : out std_logic; --  arburstm0           2   [0:1]

    AR_BUP_O2     : out std_logic; --  arburstp0           2   [0:1]
    AR_BUP_O1     : out std_logic; --  arburstp0           2   [0:1]

    AR_CHM_O4     : out std_logic; --  arcachem0           4   [0:3]
    AR_CHM_O3     : out std_logic; --  arcachem0           4   [0:3]
    AR_CHM_O2     : out std_logic; --  arcachem0           4   [0:3]
    AR_CHM_O1     : out std_logic; --  arcachem0           4   [0:3]

    AR_CHP_O4     : out std_logic; --  arcachep0           4   [0:3]
    AR_CHP_O3     : out std_logic; --  arcachep0           4   [0:3]
    AR_CHP_O2     : out std_logic; --  arcachep0           4   [0:3]
    AR_CHP_O1     : out std_logic; --  arcachep0           4   [0:3]

    AR_IDM_O4     : out std_logic; --  aridm0              4   [0:3]
    AR_IDM_O3     : out std_logic; --  aridm0              4   [0:3]
    AR_IDM_O2     : out std_logic; --  aridm0              4   [0:3]
    AR_IDM_O1     : out std_logic; --  aridm0              4   [0:3]

    AR_IDP_O4     : out std_logic; --  aridp0              4   [0:3]
    AR_IDP_O3     : out std_logic; --  aridp0              4   [0:3]
    AR_IDP_O2     : out std_logic; --  aridp0              4   [0:3]
    AR_IDP_O1     : out std_logic; --  aridp0              4   [0:3]

    AR_INM_O4     : out std_logic; --  arinnerm0           4   [0:3]
    AR_INM_O3     : out std_logic; --  arinnerm0           4   [0:3]
    AR_INM_O2     : out std_logic; --  arinnerm0           4   [0:3]
    AR_INM_O1     : out std_logic; --  arinnerm0           4   [0:3]

    AR_LEM_O4     : out std_logic; --  arlenm0             4   [0:3]
    AR_LEM_O3     : out std_logic; --  arlenm0             4   [0:3]
    AR_LEM_O2     : out std_logic; --  arlenm0             4   [0:3]
    AR_LEM_O1     : out std_logic; --  arlenm0             4   [0:3]

    AR_LEP_O4     : out std_logic; --  arlenp0             4   [0:3]
    AR_LEP_O3     : out std_logic; --  arlenp0             4   [0:3]
    AR_LEP_O2     : out std_logic; --  arlenp0             4   [0:3]
    AR_LEP_O1     : out std_logic; --  arlenp0             4   [0:3]

    AR_LKM_O2     : out std_logic; --  arlockm0            2   [0:1]
    AR_LKM_O1     : out std_logic; --  arlockm0            2   [0:1]

    AR_LKP_O2     : out std_logic; --  arlockp0            2   [0:1]
    AR_LKP_O1     : out std_logic; --  arlockp0            2   [0:1]

    AR_PRM_O3     : out std_logic; --  arprotm0            3   [0:2]
    AR_PRM_O2     : out std_logic; --  arprotm0            3   [0:2]
    AR_PRM_O1     : out std_logic; --  arprotm0            3   [0:2]

    AR_PRP_O3     : out std_logic; --  arprotp0            3   [0:2]
    AR_PRP_O2     : out std_logic; --  arprotp0            3   [0:2]
    AR_PRP_O1     : out std_logic; --  arprotp0            3   [0:2]

    AR_RDY_O      : out std_logic; --  arreadys0           1
    AR_SHM_O      : out std_logic; --  arsharem0           1

    AR_SZM_O3     : out std_logic; --  arsizem0            3   [0:2]
    AR_SZM_O2     : out std_logic; --  arsizem0            3   [0:2]
    AR_SZM_O1     : out std_logic; --  arsizem0            3   [0:2]

    AR_SZP_O3     : out std_logic; --  arsizep0            3   [0:2]
    AR_SZP_O2     : out std_logic; --  arsizep0            3   [0:2]
    AR_SZP_O1     : out std_logic; --  arsizep0            3   [0:2]

    AR_VDM_O      : out std_logic; --  arvalidm0           1
    AR_VDP_O      : out std_logic; --  arvalidp0           1

    AW_AM_O32     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O31     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O30     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O29     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O28     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O27     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O26     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O25     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O24     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O23     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O22     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O21     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O20     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O19     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O18     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O17     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O16     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O15     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O14     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O13     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O12     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O11     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O10     : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O9      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O8      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O7      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O6      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O5      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O4      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O3      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O2      : out std_logic; --  awaddrm0            32  [0:31]
    AW_AM_O1      : out std_logic; --  awaddrm0            32  [0:31]

    AW_AP_O32     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O31     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O30     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O29     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O28     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O27     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O26     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O25     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O24     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O23     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O22     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O21     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O20     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O19     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O18     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O17     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O16     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O15     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O14     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O13     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O12     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O11     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O10     : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O9      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O8      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O7      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O6      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O5      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O4      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O3      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O2      : out std_logic; --  awaddrp0            32  [0:31]
    AW_AP_O1      : out std_logic; --  awaddrp0            32  [0:31]

    AW_BUM_O2     : out std_logic; --  awburstm0           2   [0:1]
    AW_BUM_O1     : out std_logic; --  awburstm0           2   [0:1]

    AW_BUP_O2     : out std_logic; --  awburstp0           2   [0:1]
    AW_BUP_O1     : out std_logic; --  awburstp0           2   [0:1]

    AW_CHM_O4     : out std_logic; --  awcachem0           4   [0:3]
    AW_CHM_O3     : out std_logic; --  awcachem0           4   [0:3]
    AW_CHM_O2     : out std_logic; --  awcachem0           4   [0:3]
    AW_CHM_O1     : out std_logic; --  awcachem0           4   [0:3]

    AW_CHP_O4     : out std_logic; --  awcachep0           4   [0:3]
    AW_CHP_O3     : out std_logic; --  awcachep0           4   [0:3]
    AW_CHP_O2     : out std_logic; --  awcachep0           4   [0:3]
    AW_CHP_O1     : out std_logic; --  awcachep0           4   [0:3]

    AW_IDM_O4     : out std_logic; --  awidm0              4   [0:3]
    AW_IDM_O3     : out std_logic; --  awidm0              4   [0:3]
    AW_IDM_O2     : out std_logic; --  awidm0              4   [0:3]
    AW_IDM_O1     : out std_logic; --  awidm0              4   [0:3]

    AW_IDP_O4     : out std_logic; --  awidp0              4   [0:3]
    AW_IDP_O3     : out std_logic; --  awidp0              4   [0:3]
    AW_IDP_O2     : out std_logic; --  awidp0              4   [0:3]
    AW_IDP_O1     : out std_logic; --  awidp0              4   [0:3]

    AW_INM_O4     : out std_logic; --  awinnerm0           4   [0:3]
    AW_INM_O3     : out std_logic; --  awinnerm0           4   [0:3]
    AW_INM_O2     : out std_logic; --  awinnerm0           4   [0:3]
    AW_INM_O1     : out std_logic; --  awinnerm0           4   [0:3]

    AW_LEM_O4     : out std_logic; --  awlenm0             4   [0:3]
    AW_LEM_O3     : out std_logic; --  awlenm0             4   [0:3]
    AW_LEM_O2     : out std_logic; --  awlenm0             4   [0:3]
    AW_LEM_O1     : out std_logic; --  awlenm0             4   [0:3]

    AW_LEP_O4     : out std_logic; --  awlenp0             4   [0:3]
    AW_LEP_O3     : out std_logic; --  awlenp0             4   [0:3]
    AW_LEP_O2     : out std_logic; --  awlenp0             4   [0:3]
    AW_LEP_O1     : out std_logic; --  awlenp0             4   [0:3]

    AW_LKM_O2     : out std_logic; --  awlockm0            2   [0:1]
    AW_LKM_O1     : out std_logic; --  awlockm0            2   [0:1]

    AW_LKP_O2     : out std_logic; --  awlockp0            2   [0:1]
    AW_LKP_O1     : out std_logic; --  awlockp0            2   [0:1]

    AW_PRM_O3     : out std_logic; --  awprotm0            3   [0:2]
    AW_PRM_O2     : out std_logic; --  awprotm0            3   [0:2]
    AW_PRM_O1     : out std_logic; --  awprotm0            3   [0:2]

    AW_PRP_O3     : out std_logic; --  awprotp0            3   [0:2]
    AW_PRP_O2     : out std_logic; --  awprotp0            3   [0:2]
    AW_PRP_O1     : out std_logic; --  awprotp0            3   [0:2]

    AW_RDY_O      : out std_logic; --  awreadys0           1
    AW_SHM_O      : out std_logic; --  awsharem0           1

    AW_SZM_O3     : out std_logic; --  awsizem0            3   [0:2]
    AW_SZM_O2     : out std_logic; --  awsizem0            3   [0:2]
    AW_SZM_O1     : out std_logic; --  awsizem0            3   [0:2]

    AW_SZP_O3     : out std_logic; --  awsizep0            3   [0:2]
    AW_SZP_O2     : out std_logic; --  awsizep0            3   [0:2]
    AW_SZP_O1     : out std_logic; --  awsizep0            3   [0:2]

    AW_VDM_O      : out std_logic; --  awvalidm0           1
    AW_VDP_O      : out std_logic; --  awvalidp0           1

    B_IDS_O8      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O7      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O6      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O5      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O4      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O3      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O2      : out std_logic; --  bids0               8   [0:7]
    B_IDS_O1      : out std_logic; --  bids0               8   [0:7]

    B_RDYM_O      : out std_logic; --  breadym0            1
    B_RDYP_O      : out std_logic; --  breadyp0            1

    B_RSP_O2      : out std_logic; --  bresps0             2   [0:1]
    B_RSP_O1      : out std_logic; --  bresps0             2   [0:1]

    B_VD_O        : out std_logic; --  bvalids0            1

--    CAL_O5        : out std_logic; --  calibration         5   [0:4]
--    CAL_O4        : out std_logic; --  calibration         5   [0:4]
--    CAL_O3        : out std_logic; --  calibration         5   [0:4]
--    CAL_O2        : out std_logic; --  calibration         5   [0:4]
--    CAL_O1        : out std_logic; --  calibration         5   [0:4]

    CDB_PW_O      : out std_logic; --  cdbgpwrupreq        1
    CDB_RS_O      : out std_logic; --  cdbgrstreq          1
--    CK_DR_O       : out std_logic; --  clock_dr            1
    COM_RX_O      : out std_logic; --  commrx0             1
    COM_TX_O      : out std_logic; --  commtx0             1
    CS_PW_O       : out std_logic; --  csyspwrupreq        1
    DB_ACK_O      : out std_logic; --  dbgack0             1
    DB_NPD_O      : out std_logic; --  dbgnopwrdwn         1
    DB_RS_O       : out std_logic; --  dbgrstreq0          1

    DFTS_O8       : out std_logic; --  dftso               8   [0:7]
    DFTS_O7       : out std_logic; --  dftso               8   [0:7]
    DFTS_O6       : out std_logic; --  dftso               8   [0:7]
    DFTS_O5       : out std_logic; --  dftso               8   [0:7]
    DFTS_O4       : out std_logic; --  dftso               8   [0:7]
    DFTS_O3       : out std_logic; --  dftso               8   [0:7]
    DFTS_O2       : out std_logic; --  dftso               8   [0:7]
    DFTS_O1       : out std_logic; --  dftso               8   [0:7]

    ET_ASC_O8     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O7     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O6     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O5     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O4     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O3     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O2     : out std_logic; --  etmasicctl0         8   [0:7]
    ET_ASC_O1     : out std_logic; --  etmasicctl0         8   [0:7]

    ET_E_O        : out std_logic; --  etmen0              1

    ET_EXT_O2     : out std_logic; --  etmextout0          2   [0:1]
    ET_EXT_O1     : out std_logic; --  etmextout0          2   [0:1]

    EVENT_O       : out std_logic; --  evento0             1
    FP_DZC_O      : out std_logic; --  fpdzc0              1
    FP_IDC_O      : out std_logic; --  fpidc0              1
    FP_IOC_O      : out std_logic; --  fpioc0              1
    FP_IXC_O      : out std_logic; --  fpixc0              1
    FP_OFC_O      : out std_logic; --  fpofc0              1
    FP_UFC_O      : out std_logic; --  fpufc0              1
    JTAG_O        : out std_logic; --  jtagnsw             1
--    LBK_E_O       : out std_logic; --  loopback_en         1
--    LBK_MX_O      : out std_logic; --  loopback_mux        1

--    MODE1_O2      : out std_logic; --  mode1               3   [0:2]
--    MODE1_O1      : out std_logic; --  mode1               3   [0:2]

--    MODE2_O2      : out std_logic; --  mode2               3   [0:2]
--    MODE2_O1      : out std_logic; --  mode2               3   [0:2]

--    MODE3_O2      : out std_logic; --  mode3               3   [0:2]
--    MODE3_O1      : out std_logic; --  mode3               3   [0:2]

    N_CKST_O      : out std_logic; --  nclkstopped0        1
    N_PMU_O       : out std_logic; --  npmuirq0            1
    N_TDO_O       : out std_logic; --  ntdoen              1
    N_VFIQ_O      : out std_logic; --  nvalfiq0            1
    N_VIRQ_O      : out std_logic; --  nvalirq0            1
    N_VRST_O      : out std_logic; --  nvalreset0          1
    N_EPST_O      : out std_logic; --  nwfepipestopped0    1
    N_IPST_O      : out std_logic; --  nwfipipestopped0    1

    P_RD_O32      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O31      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O30      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O29      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O28      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O27      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O26      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O25      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O24      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O23      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O22      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O21      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O20      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O19      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O18      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O17      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O16      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O15      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O14      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O13      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O12      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O11      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O10      : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O9       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O8       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O7       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O6       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O5       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O4       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O3       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O2       : out std_logic; --  prdatasys           32  [0:31]
    P_RD_O1       : out std_logic; --  prdatasys           32  [0:31]

    P_RDY_O       : out std_logic; --  preadysys           1
    P_VER_O       : out std_logic; --  pslverrsys          1

    RD_O64        : out std_logic; --  rdatas0             64  [0:63]
    RD_O63        : out std_logic; --  rdatas0             64  [0:63]
    RD_O62        : out std_logic; --  rdatas0             64  [0:63]
    RD_O61        : out std_logic; --  rdatas0             64  [0:63]
    RD_O60        : out std_logic; --  rdatas0             64  [0:63]
    RD_O59        : out std_logic; --  rdatas0             64  [0:63]
    RD_O58        : out std_logic; --  rdatas0             64  [0:63]
    RD_O57        : out std_logic; --  rdatas0             64  [0:63]
    RD_O56        : out std_logic; --  rdatas0             64  [0:63]
    RD_O55        : out std_logic; --  rdatas0             64  [0:63]
    RD_O54        : out std_logic; --  rdatas0             64  [0:63]
    RD_O53        : out std_logic; --  rdatas0             64  [0:63]
    RD_O52        : out std_logic; --  rdatas0             64  [0:63]
    RD_O51        : out std_logic; --  rdatas0             64  [0:63]
    RD_O50        : out std_logic; --  rdatas0             64  [0:63]
    RD_O49        : out std_logic; --  rdatas0             64  [0:63]
    RD_O48        : out std_logic; --  rdatas0             64  [0:63]
    RD_O47        : out std_logic; --  rdatas0             64  [0:63]
    RD_O46        : out std_logic; --  rdatas0             64  [0:63]
    RD_O45        : out std_logic; --  rdatas0             64  [0:63]
    RD_O44        : out std_logic; --  rdatas0             64  [0:63]
    RD_O43        : out std_logic; --  rdatas0             64  [0:63]
    RD_O42        : out std_logic; --  rdatas0             64  [0:63]
    RD_O41        : out std_logic; --  rdatas0             64  [0:63]
    RD_O40        : out std_logic; --  rdatas0             64  [0:63]
    RD_O39        : out std_logic; --  rdatas0             64  [0:63]
    RD_O38        : out std_logic; --  rdatas0             64  [0:63]
    RD_O37        : out std_logic; --  rdatas0             64  [0:63]
    RD_O36        : out std_logic; --  rdatas0             64  [0:63]
    RD_O35        : out std_logic; --  rdatas0             64  [0:63]
    RD_O34        : out std_logic; --  rdatas0             64  [0:63]
    RD_O33        : out std_logic; --  rdatas0             64  [0:63]
    RD_O32        : out std_logic; --  rdatas0             64  [0:63]
    RD_O31        : out std_logic; --  rdatas0             64  [0:63]
    RD_O30        : out std_logic; --  rdatas0             64  [0:63]
    RD_O29        : out std_logic; --  rdatas0             64  [0:63]
    RD_O28        : out std_logic; --  rdatas0             64  [0:63]
    RD_O27        : out std_logic; --  rdatas0             64  [0:63]
    RD_O26        : out std_logic; --  rdatas0             64  [0:63]
    RD_O25        : out std_logic; --  rdatas0             64  [0:63]
    RD_O24        : out std_logic; --  rdatas0             64  [0:63]
    RD_O23        : out std_logic; --  rdatas0             64  [0:63]
    RD_O22        : out std_logic; --  rdatas0             64  [0:63]
    RD_O21        : out std_logic; --  rdatas0             64  [0:63]
    RD_O20        : out std_logic; --  rdatas0             64  [0:63]
    RD_O19        : out std_logic; --  rdatas0             64  [0:63]
    RD_O18        : out std_logic; --  rdatas0             64  [0:63]
    RD_O17        : out std_logic; --  rdatas0             64  [0:63]
    RD_O16        : out std_logic; --  rdatas0             64  [0:63]
    RD_O15        : out std_logic; --  rdatas0             64  [0:63]
    RD_O14        : out std_logic; --  rdatas0             64  [0:63]
    RD_O13        : out std_logic; --  rdatas0             64  [0:63]
    RD_O12        : out std_logic; --  rdatas0             64  [0:63]
    RD_O11        : out std_logic; --  rdatas0             64  [0:63]
    RD_O10        : out std_logic; --  rdatas0             64  [0:63]
    RD_O9         : out std_logic; --  rdatas0             64  [0:63]
    RD_O8         : out std_logic; --  rdatas0             64  [0:63]
    RD_O7         : out std_logic; --  rdatas0             64  [0:63]
    RD_O6         : out std_logic; --  rdatas0             64  [0:63]
    RD_O5         : out std_logic; --  rdatas0             64  [0:63]
    RD_O4         : out std_logic; --  rdatas0             64  [0:63]
    RD_O3         : out std_logic; --  rdatas0             64  [0:63]
    RD_O2         : out std_logic; --  rdatas0             64  [0:63]
    RD_O1         : out std_logic; --  rdatas0             64  [0:63]

--    RDY_O3        : out std_logic; --  ready               3   [0:2]
--    RDY_O2        : out std_logic; --  ready               3   [0:2]
--    RDY_O1        : out std_logic; --  ready               3   [0:2]

    R_IDS_O8      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O7      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O6      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O5      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O4      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O3      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O2      : out std_logic; --  rids0               8   [0:7]
    R_IDS_O1      : out std_logic; --  rids0               8   [0:7]

    R_LST_O       : out std_logic; --  rlasts0             1
    R_RDYM_O      : out std_logic; --  rreadym0            1
    R_RDYP_O      : out std_logic; --  rreadyp0            1

    R_RSP_O2      : out std_logic; --  rresps0             2   [0:1]
    R_RSP_O1      : out std_logic; --  rresps0             2   [0:1]

    R_VD_O        : out std_logic; --  rvalids0            1
--    SCAN_E_O      : out std_logic; --  scan_en             1
--    SHF_DR_O      : out std_logic; --  shift_dr            1
--    SHOUT_O       : out std_logic; --  shout               1
    SWDO_O        : out std_logic; --  swdo                1
    SWDO_E_O      : out std_logic; --  swdoen              1
    TDO_O         : out std_logic; --  tdo                 1
--    TEST_E_O      : out std_logic; --  test_en             1
    T_CK_O        : out std_logic; --  traceclk            1
    T_CTL_O       : out std_logic; --  tracectl            1

    T_DATA_O32    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O31    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O30    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O29    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O28    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O27    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O26    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O25    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O24    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O23    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O22    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O21    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O20    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O19    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O18    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O17    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O16    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O15    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O14    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O13    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O12    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O11    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O10    : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O9     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O8     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O7     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O6     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O5     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O4     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O3     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O2     : out std_logic; --  tracedata           32  [0:31]
    T_DATA_O1     : out std_logic; --  tracedata           32  [0:31]

--    UPD_DR_O      : out std_logic; --  update_dr           1

    W_DM_O64      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O63      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O62      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O61      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O60      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O59      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O58      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O57      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O56      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O55      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O54      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O53      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O52      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O51      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O50      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O49      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O48      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O47      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O46      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O45      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O44      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O43      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O42      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O41      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O40      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O39      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O38      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O37      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O36      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O35      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O34      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O33      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O32      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O31      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O30      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O29      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O28      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O27      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O26      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O25      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O24      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O23      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O22      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O21      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O20      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O19      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O18      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O17      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O16      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O15      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O14      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O13      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O12      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O11      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O10      : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O9       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O8       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O7       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O6       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O5       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O4       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O3       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O2       : out std_logic; --  wdatam0             64  [0:63]
    W_DM_O1       : out std_logic; --  wdatam0             64  [0:63]

    W_DP_O32      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O31      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O30      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O29      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O28      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O27      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O26      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O25      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O24      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O23      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O22      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O21      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O20      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O19      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O18      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O17      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O16      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O15      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O14      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O13      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O12      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O11      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O10      : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O9       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O8       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O7       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O6       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O5       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O4       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O3       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O2       : out std_logic; --  wdatap0             32  [0:31]
    W_DP_O1       : out std_logic; --  wdatap0             32  [0:31]

    W_IDM_O4      : out std_logic; --  widm0               4   [0:3]
    W_IDM_O3      : out std_logic; --  widm0               4   [0:3]
    W_IDM_O2      : out std_logic; --  widm0               4   [0:3]
    W_IDM_O1      : out std_logic; --  widm0               4   [0:3]

    W_IDP_O4      : out std_logic; --  widp0               4   [0:3]
    W_IDP_O3      : out std_logic; --  widp0               4   [0:3]
    W_IDP_O2      : out std_logic; --  widp0               4   [0:3]
    W_IDP_O1      : out std_logic; --  widp0               4   [0:3]

    W_LSTM_O      : out std_logic; --  wlastm0             1
    W_LSTP_O      : out std_logic; --  wlastp0             1
    W_RDY_O       : out std_logic; --  wreadys0            1

    W_SBM_O8      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O7      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O6      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O5      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O4      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O3      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O2      : out std_logic; --  wstrbm0             8   [0:7]
    W_SBM_O1      : out std_logic; --  wstrbm0             8   [0:7]

    W_SBP_O4      : out std_logic; --  wstrbp0             4   [0:3]
    W_SBP_O3      : out std_logic; --  wstrbp0             4   [0:3]
    W_SBP_O2      : out std_logic; --  wstrbp0             4   [0:3]
    W_SBP_O1      : out std_logic; --  wstrbp0             4   [0:3]

    W_VDM_O       : out std_logic; --  wvalidm0            1
    W_VDP_O       : out std_logic  --  wvalidp0            1
);
end NX_R5_L;

-- =================================================================================================
--   NX_R5_L_WRAP definition                                                            2019/04/09
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_R5_L_WRAP is
port (
            ------------------------------------------------------------------------
            -- CORTEXR5 PRIMARY INPUTS AND OUTPUTS
            ------------------------------------------------------------------------  
            ------------------------------------------------------------------------
            -- Global
            ------------------------------------------------------------------------
            CLKIN                  : in std_logic;
            nRESET0                : in std_logic;
            nSYSPORESET            : in std_logic;
            nCPUHALT0              : in std_logic;
            DBGNOCLKSTOP           : in std_logic;
            nCLKSTOPPED0           : out std_logic;
            nWFEPIPESTOPPED0       : out std_logic;
            nWFIPIPESTOPPED0       : out std_logic;
            EVENTI0                : in std_logic;
            EVENTO0                : out std_logic;
            ------------------------------------------------------------------------
            -- Configuration signals
            ------------------------------------------------------------------------
            VINITHI0               : in std_logic;        
            CFGEE                  : in std_logic;        
            CFGIE                  : in std_logic;        
            INITRAMA0              : in std_logic;        
            LOCZRAMA0              : in std_logic;        
            TEINIT                 : in std_logic;        
            CFGNMFI0               : in std_logic;        
            PARECCENRAM0           : in std_logic;        
            PARITYLEVEL            : in std_logic;        
            ERRENRAM0              : in std_logic;        
            GROUPID                : in std_logic_vector(3 downto 0);        
            INITPPX0               : in std_logic;        
            PPXBASE0               : in std_logic_vector(19 downto 0);        
            PPXSIZE0               : in std_logic_vector(4 downto 0);        
            PPVBASE0               : in std_logic_vector(19 downto 0);        
            PPVSIZE0               : in std_logic_vector(4 downto 0);        
            ------------------------------------------------------------------------
            -- Interrupt signals
            ------------------------------------------------------------------------
            nFIQ0          : in std_logic;        
            nIRQ0          : in std_logic;        
            nPMUIRQ0       : out std_logic;        
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Master Port
            ------------------------------------------------------------------------
            ACLKENM0       : in std_logic;       
            -- Write Address Channel
            AWADDRM0       : out std_logic_vector(31 downto 0);        
            AWBURSTM0      : out std_logic_vector(1 downto 0);        
            AWCACHEM0      : out std_logic_vector(3 downto 0);        
            AWIDM0         : out std_logic_vector(3 downto 0);        
            AWLENM0        : out std_logic_vector(3 downto 0);        
            AWLOCKM0       : out std_logic_vector(1 downto 0);        
            AWPROTM0       : out std_logic_vector(2 downto 0);        
            AWREADYM0      : in std_logic;        
            AWSIZEM0       : out std_logic_vector(2 downto 0);       
            AWINNERM0      : out std_logic_vector(3 downto 0);       
            AWSHAREM0      : out std_logic;       
            AWVALIDM0      : out std_logic;       
            -- Write Data Channel
            WDATAM0        : out std_logic_vector(63 downto 0);       
            WIDM0          : out std_logic_vector(3 downto 0);       
            WLASTM0        : out std_logic;       
            WREADYM0       : in std_logic;       
            WSTRBM0        : out std_logic_vector(7 downto 0);       
            WVALIDM0       : out std_logic;       
            -- Write response channel
            BIDM0           : in std_logic_vector(3 downto 0);       
            BREADYM0        : out std_logic;       
            BRESPM0         : in std_logic_vector(1 downto 0);       
            BVALIDM0        : in std_logic;       
            -- Read Address Channel
            ARADDRM0    : out std_logic_vector(31 downto 0);          
            ARBURSTM0   : out std_logic_vector(1 downto 0);          
            ARCACHEM0   : out std_logic_vector(3 downto 0);          
            ARIDM0      : out std_logic_vector(3 downto 0);          
            ARLENM0     : out std_logic_vector(3 downto 0);          
            ARLOCKM0    : out std_logic_vector(1 downto 0);          
            ARPROTM0    : out std_logic_vector(2 downto 0);          
            ARREADYM0   : in std_logic;          
            ARSIZEM0    : out std_logic_vector(2 downto 0);           
            ARINNERM0   : out std_logic_vector(3 downto 0);           
            ARSHAREM0   : out std_logic;           
            ARVALIDM0   : out std_logic;           
            -- Read Data Channel
            RDATAM0     : in std_logic_vector(63 downto 0);           
            RIDM0       : in std_logic_vector(3 downto 0);           
            RLASTM0     : in std_logic;           
            RREADYM0    : out std_logic;           
            RRESPM0     : in std_logic_vector(1 downto 0);           
            RVALIDM0    : in std_logic;           
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Slave Port
            ------------------------------------------------------------------------
            ACLKENS0    : in std_logic;           
            -- Write Address Channel
            AWADDRS0    : in std_logic_vector(31 downto 0);           
            AWBURSTS0   : in std_logic_vector(1 downto 0);           
            AWCACHES0   : in std_logic_vector(3 downto 0);           

            AWIDS0      : in std_logic_vector(7 downto 0);           
            AWLENS0     : in std_logic_vector(3 downto 0);           
            AWLOCKS0    : in std_logic_vector(1 downto 0);           
            AWPROTS0    : in std_logic_vector(2 downto 0);           
            AWREADYS0   : out std_logic;          
            AWSIZES0    : in std_logic_vector(2 downto 0);           
            AWVALIDS0   : in std_logic;           
            -- Write Data Channel
            WDATAS0     : in std_logic_vector(63 downto 0);           
            WIDS0       : in std_logic_vector(7 downto 0);           
            WLASTS0     : in std_logic;           
            WREADYS0    : out std_logic;           
            WSTRBS0     : in std_logic_vector(7 downto 0);          
            WVALIDS0    : in std_logic;           
            -- Write response channel
            BIDS0       : out std_logic_vector(7 downto 0);           
            BREADYS0    : in std_logic;           
            BRESPS0     : out std_logic_vector(1 downto 0);           
            BVALIDS0    : out std_logic;           
            -- Read Address Channel
            ARADDRS0    : in std_logic_vector(31 downto 0);           
            ARBURSTS0   : in std_logic_vector(1 downto 0);           
            ARCACHES0   : in std_logic_vector(3 downto 0);           
            ARIDS0      : in std_logic_vector(7 downto 0);           
            ARLENS0     : in std_logic_vector(3 downto 0);           
            ARLOCKS0    : in std_logic_vector(1 downto 0);           
            ARPROTS0    : in std_logic_vector(2 downto 0);           
            ARREADYS0   : out std_logic;           
            ARSIZES0    : in std_logic_vector(2 downto 0);           

            ARVALIDS0   : in std_logic;           
            -- Read Data Channel
            RDATAS0     : out std_logic_vector(63 downto 0);           
            RIDS0       : out std_logic_vector(7 downto 0);           
            RLASTS0     : out std_logic;           
            RREADYS0    : in std_logic;           
            RRESPS0     : out std_logic_vector(1 downto 0);           
            RVALIDS0    : out std_logic;           
            ------------------------------------------------------------------------
            -- L2 interface signals - AXI Peripheral Port
            ------------------------------------------------------------------------
            ACLKENP0     : in std_logic;          
            -- Write Address Channel
            AWIDP0       : out std_logic_vector(3 downto 0);          
            AWADDRP0     : out std_logic_vector(31 downto 0);          
            AWLENP0      : out std_logic_vector(3 downto 0);          
            AWSIZEP0     : out std_logic_vector(2 downto 0);          
            AWBURSTP0    : out std_logic_vector(1 downto 0);          
            AWLOCKP0     : out std_logic_vector(1 downto 0);          
            AWCACHEP0    : out std_logic_vector(3 downto 0);          
            AWPROTP0     : out std_logic_vector(2 downto 0);          
            AWVALIDP0    : out std_logic;          
            AWREADYP0    : in std_logic;          
            -- Write Data Channel
            WIDP0        : out std_logic_vector(3 downto 0);          
            WDATAP0      : out std_logic_vector(31 downto 0);          
            WSTRBP0      : out std_logic_vector(3 downto 0);          
            WLASTP0      : out std_logic;          
            WVALIDP0     : out std_logic;          
            WREADYP0     : in std_logic;          
            -- Write response channel
            BIDP0        : in std_logic_vector(3 downto 0);          
            BRESPP0      : in std_logic_vector(1 downto 0);          
            BVALIDP0     : in std_logic;          
            BREADYP0     : out std_logic;          
            -- Read Address Channel
            ARIDP0       : out std_logic_vector (3 downto 0);          
            ARADDRP0     : out std_logic_vector (31 downto 0);          
            ARLENP0      : out std_logic_vector (3 downto 0);          
            ARSIZEP0     : out std_logic_vector (2 downto 0);          
            ARBURSTP0    : out std_logic_vector (1 downto 0);          
            ARLOCKP0     : out std_logic_vector (1 downto 0);          
            ARCACHEP0    : out std_logic_vector (3 downto 0);          
            ARPROTP0     : out std_logic_vector (2 downto 0);          
            ARVALIDP0    : out std_logic;          
            ARREADYP0    : in std_logic;          
            -- Reainata Channel
            RIDP0        : in std_logic_vector(3 downto 0);          
            RDATAP0      : in std_logic_vector(31 downto 0);          
            RRESPP0      : in std_logic_vector(1 downto 0);          
            RLASTP0      : in std_logic;          
            RVALIDP0     : in std_logic;          
            RREADYP0     : out std_logic;          
       
            -- Debug Miscellaneous
            DBGEN0       : in std_logic;          
            NIDEN0       : in std_logic;          
            EDBGRQ0      : in std_logic;          
            DBGACK0      : out std_logic;          
            DBGRSTREQ0   : out std_logic;          

            COMMRX0      : out std_logic;          
            COMMTX0      : out std_logic;          

            DBGNOPWRDWN    : out std_logic;        
            DBGROMADDR     : in std_logic_vector(19 downto 0);        
            DBGROMADDRV    : in std_logic;        
            DBGSELFADDR0   : in std_logic_vector(19 downto 0);        
            DBGSELFADDRV0  : in std_logic;        
            ------------------------------------------------------------------------
            -- ETM Interface
            ------------------------------------------------------------------------
            nETMPORESET    : in std_logic;        
            ETMASICCTL0    : out std_logic_vector(7 downto 0);        
            ETMEN0         : out std_logic;        
            ETMEXTOUT0     : out std_logic_vector(1 downto 0);        
            ------------------------------------------------------------------------
            -- Validation
            ------------------------------------------------------------------------
            nVALIRQ0        : out std_logic;       
            nVALFIQ0        : out std_logic;       
            nVALRESET0      : out std_logic;       
       
            ------------------------------------------------------------------------
            -- FPU
            ------------------------------------------------------------------------
           FPIXC0           : out std_logic;      
           FPOFC0           : out std_logic;      
           FPUFC0           : out std_logic;      
           FPIOC0           : out std_logic;      
           FPDZC0           : out std_logic;      
           FPIDC0           : out std_logic;      
            ------------------------------------------------------------------------
            -- Coresight TPIU-Lite
            ------------------------------------------------------------------------
            ------------------------------------------------------------------------
            -- ATB Port
            ------------------------------------------------------------------------
            ATRESETn   : in std_logic;            
            ------------------------------------------------------------------------
            -- Trace Out Port
            ------------------------------------------------------------------------
            TRACECLK     : out std_logic;          
            TRACEDATA    : out std_logic_vector(31 downto 0);          
            TRACECTL     : out std_logic;          
            ------------------------------------------------------------------------
            -- Coresight DAP-Lite
            ------------------------------------------------------------------------
            ------------------------------------------------------------------------
            -- CoreSight DAP Ports
            ------------------------------------------------------------------------    
            PCLKSYS           : in std_logic;     
            PCLKENSYS         : in std_logic;     
            PRESETSYSn        : in std_logic;     
            PADDRSYS          : in std_logic_vector(28 downto 0);     
            PENABLESYS        : in std_logic;     
            PRDATASYS         : out std_logic_vector(31 downto 0);     
            PREADYSYS         : out std_logic;     
            PSELSYS           : in std_logic;     
            PSLVERRSYS        : out std_logic;     
            PWDATASYS         : in std_logic_vector(31 downto 0);     
            PWRITESYS         : in std_logic;     
       
            CDBGPWRUPACK       : in std_logic;    
            CDBGPWRUPREQ       : out std_logic;    
            CDBGRSTACK         : in std_logic;    
            CDBGRSTREQ         : out std_logic;    
            CSYSPWRUPACK       : in std_logic;    
            CSYSPWRUPREQ       : out std_logic;    
            DEVICEEN           : in std_logic;    
            JTAGNSW            : out std_logic;    
            nPOTRST            : in std_logic;    
            nTDOEN             : out std_logic;    
            nTRST              : in std_logic;    
            SWCLKTCK           : in std_logic;    
            SWDITMS            : in std_logic;    
            SWDO               : out std_logic;    
            SWDOEN             : out std_logic;    
            TDI                : in std_logic;    
            TDO                : out std_logic    

);
end NX_R5_L_WRAP;

architecture NX_RTL of NX_R5_L_WRAP is
begin

    inst_NX_R : NX_R5_L
    port map (
	-- Inputs
	  A_CKEM_I      =>  ACLKENM0
	, A_CKEP_I      =>  ACLKENP0
	, A_CKES_I      =>  ACLKENS0

	, AR_A_I32      =>  ARADDRS0(31)
	, AR_A_I31      =>  ARADDRS0(30)
	, AR_A_I30      =>  ARADDRS0(29)
	, AR_A_I29      =>  ARADDRS0(28)
	, AR_A_I28      =>  ARADDRS0(27)
	, AR_A_I27      =>  ARADDRS0(26)
	, AR_A_I26      =>  ARADDRS0(25)
	, AR_A_I25      =>  ARADDRS0(24)
	, AR_A_I24      =>  ARADDRS0(23)
	, AR_A_I23      =>  ARADDRS0(22)
	, AR_A_I22      =>  ARADDRS0(21)
	, AR_A_I21      =>  ARADDRS0(20)
	, AR_A_I20      =>  ARADDRS0(19)
	, AR_A_I19      =>  ARADDRS0(18)
	, AR_A_I18      =>  ARADDRS0(17)
	, AR_A_I17      =>  ARADDRS0(16)
	, AR_A_I16      =>  ARADDRS0(15)
	, AR_A_I15      =>  ARADDRS0(14)
	, AR_A_I14      =>  ARADDRS0(13)
	, AR_A_I13      =>  ARADDRS0(12)
	, AR_A_I12      =>  ARADDRS0(11)
	, AR_A_I11      =>  ARADDRS0(10)
	, AR_A_I10      =>  ARADDRS0(9)
	, AR_A_I9       =>  ARADDRS0(8)
	, AR_A_I8       =>  ARADDRS0(7)
	, AR_A_I7       =>  ARADDRS0(6)
	, AR_A_I6       =>  ARADDRS0(5)
	, AR_A_I5       =>  ARADDRS0(4)
	, AR_A_I4       =>  ARADDRS0(3)
	, AR_A_I3       =>  ARADDRS0(2)
	, AR_A_I2       =>  ARADDRS0(1)
	, AR_A_I1       =>  ARADDRS0(0)

	, AR_BU_I2      =>  ARBURSTS0(1)
	, AR_BU_I1      =>  ARBURSTS0(0)

	, AR_CH_I4      =>  ARCACHES0(3)
	, AR_CH_I3      =>  ARCACHES0(2)
	, AR_CH_I2      =>  ARCACHES0(1)
	, AR_CH_I1      =>  ARCACHES0(0)

	, AR_IDS_I8     =>  ARIDS0(7)
	, AR_IDS_I7     =>  ARIDS0(6)
	, AR_IDS_I6     =>  ARIDS0(5)
	, AR_IDS_I5     =>  ARIDS0(4)
	, AR_IDS_I4     =>  ARIDS0(3)
	, AR_IDS_I3     =>  ARIDS0(2)
	, AR_IDS_I2     =>  ARIDS0(1)
	, AR_IDS_I1     =>  ARIDS0(0)

	, AR_LE_I4      =>  ARLENS0(3)
	, AR_LE_I3      =>  ARLENS0(2)
	, AR_LE_I2      =>  ARLENS0(1)
	, AR_LE_I1      =>  ARLENS0(0)

	, AR_LK_I2      =>  ARLOCKS0(1)
	, AR_LK_I1      =>  ARLOCKS0(0)

	, AR_PR_I3      =>  ARPROTS0(2)
	, AR_PR_I2      =>  ARPROTS0(1)
	, AR_PR_I1      =>  ARPROTS0(0)

	, AR_RYM_I      =>  ARREADYM0
	, AR_RYP_I      =>  ARREADYP0

	, AR_SZ_I3      =>  ARSIZES0(2)
	, AR_SZ_I2      =>  ARSIZES0(1)
	, AR_SZ_I1      =>  ARSIZES0(0)

	, AR_VD_I       =>  ARVALIDS0
	, AT_RS_I       =>  ATRESETn

	, AW_A_I32      =>  AWADDRS0(31)
	, AW_A_I31      =>  AWADDRS0(30)
	, AW_A_I30      =>  AWADDRS0(29)
	, AW_A_I29      =>  AWADDRS0(28)
	, AW_A_I28      =>  AWADDRS0(27)
	, AW_A_I27      =>  AWADDRS0(26)
	, AW_A_I26      =>  AWADDRS0(25)
	, AW_A_I25      =>  AWADDRS0(24)
	, AW_A_I24      =>  AWADDRS0(23)
	, AW_A_I23      =>  AWADDRS0(22)
	, AW_A_I22      =>  AWADDRS0(21)
	, AW_A_I21      =>  AWADDRS0(20)
	, AW_A_I20      =>  AWADDRS0(19)
	, AW_A_I19      =>  AWADDRS0(18)
	, AW_A_I18      =>  AWADDRS0(17)
	, AW_A_I17      =>  AWADDRS0(16)
	, AW_A_I16      =>  AWADDRS0(15)
	, AW_A_I15      =>  AWADDRS0(14)
	, AW_A_I14      =>  AWADDRS0(13)
	, AW_A_I13      =>  AWADDRS0(12)
	, AW_A_I12      =>  AWADDRS0(11)
	, AW_A_I11      =>  AWADDRS0(10)
	, AW_A_I10      =>  AWADDRS0(9)
	, AW_A_I9       =>  AWADDRS0(8)
	, AW_A_I8       =>  AWADDRS0(7)
	, AW_A_I7       =>  AWADDRS0(6)
	, AW_A_I6       =>  AWADDRS0(5)
	, AW_A_I5       =>  AWADDRS0(4)
	, AW_A_I4       =>  AWADDRS0(3)
	, AW_A_I3       =>  AWADDRS0(2)
	, AW_A_I2       =>  AWADDRS0(1)
	, AW_A_I1       =>  AWADDRS0(0)

	, AW_BU_I2      =>  AWBURSTS0(1)
	, AW_BU_I1      =>  AWBURSTS0(0)

	, AW_CH_I4      =>  AWCACHES0(3)
	, AW_CH_I3      =>  AWCACHES0(2)
	, AW_CH_I2      =>  AWCACHES0(1)
	, AW_CH_I1      =>  AWCACHES0(0)

	, AW_IDS_I8     =>  AWIDS0(7)
	, AW_IDS_I7     =>  AWIDS0(6)
	, AW_IDS_I6     =>  AWIDS0(5)
	, AW_IDS_I5     =>  AWIDS0(4)
	, AW_IDS_I4     =>  AWIDS0(3)
	, AW_IDS_I3     =>  AWIDS0(2)
	, AW_IDS_I2     =>  AWIDS0(1)
	, AW_IDS_I1     =>  AWIDS0(0)

	, AW_LE_I4      =>  AWLENS0(3)
	, AW_LE_I3      =>  AWLENS0(2)
	, AW_LE_I2      =>  AWLENS0(1)
	, AW_LE_I1      =>  AWLENS0(0)

	, AW_LK_I2      =>  AWLOCKS0(1)
	, AW_LK_I1      =>  AWLOCKS0(0)

	, AW_PR_I3      =>  AWPROTS0(2)
	, AW_PR_I2      =>  AWPROTS0(1)
	, AW_PR_I1      =>  AWPROTS0(0)

	, AW_RYM_I      =>  AWREADYM0
	, AW_RYP_I      =>  AWREADYP0

	, AW_SZ_I3      =>  AWSIZES0(2)
	, AW_SZ_I2      =>  AWSIZES0(1)
	, AW_SZ_I1      =>  AWSIZES0(0)

	, AW_VD_I       =>  AWVALIDS0

	, B_IDM_I4      =>  BIDM0(3)
	, B_IDM_I3      =>  BIDM0(2)
	, B_IDM_I2      =>  BIDM0(1)
	, B_IDM_I1      =>  BIDM0(0)

	, B_IDP_I4      =>  BIDP0(3)
	, B_IDP_I3      =>  BIDP0(2)
	, B_IDP_I2      =>  BIDP0(1)
	, B_IDP_I1      =>  BIDP0(0)

	, B_RDY_I       =>  BREADYS0

	, B_RSPM_I2     =>  BRESPM0(1)
	, B_RSPM_I1     =>  BRESPM0(0)

	, B_RSPP_I2     =>  BRESPP0(1)
	, B_RSPP_I1     =>  BRESPP0(0)

	, B_VDM_I       =>  BVALIDM0
	, B_VDP_I       =>  BVALIDP0

--	, CAL_I5        =>  CAL_I(4)
--	, CAL_I4        =>  CAL_I(3)
--	, CAL_I3        =>  CAL_I(2)
--	, CAL_I2        =>  CAL_I(1)
--	, CAL_I1        =>  CAL_I(0)

	, CDB_PW_I      =>  CDBGPWRUPACK
	, CDB_RS_I      =>  CDBGRSTACK
	, CFG_EE_I      =>  CFGEE
	, CFG_IE_I      =>  CFGIE
	, CFG_NM_I      =>  CFGNMFI0
	, CK_I          =>  CLKIN
--	, CK_DR_I       =>  CK_DR_I
	, CS_PW_I       =>  CSYSPWRUPACK
	, DB_E_I        =>  DBGEN0
	, DB_NCK_I      =>  DBGNOCLKSTOP

	, DB_RA_I20     =>  DBGROMADDR(19)
	, DB_RA_I19     =>  DBGROMADDR(18)
	, DB_RA_I18     =>  DBGROMADDR(17)
	, DB_RA_I17     =>  DBGROMADDR(16)
	, DB_RA_I16     =>  DBGROMADDR(15)
	, DB_RA_I15     =>  DBGROMADDR(14)
	, DB_RA_I14     =>  DBGROMADDR(13)
	, DB_RA_I13     =>  DBGROMADDR(12)
	, DB_RA_I12     =>  DBGROMADDR(11)
	, DB_RA_I11     =>  DBGROMADDR(10)
	, DB_RA_I10     =>  DBGROMADDR(9)
	, DB_RA_I9      =>  DBGROMADDR(8)
	, DB_RA_I8      =>  DBGROMADDR(7)
	, DB_RA_I7      =>  DBGROMADDR(6)
	, DB_RA_I6      =>  DBGROMADDR(5)
	, DB_RA_I5      =>  DBGROMADDR(4)
	, DB_RA_I4      =>  DBGROMADDR(3)
	, DB_RA_I3      =>  DBGROMADDR(2)
	, DB_RA_I2      =>  DBGROMADDR(1)
	, DB_RA_I1      =>  DBGROMADDR(0)

	, DB_RAV_I      =>  DBGROMADDRV

	, DB_SA_I20     =>  DBGSELFADDR0(19)
	, DB_SA_I19     =>  DBGSELFADDR0(18)
	, DB_SA_I18     =>  DBGSELFADDR0(17)
	, DB_SA_I17     =>  DBGSELFADDR0(16)
	, DB_SA_I16     =>  DBGSELFADDR0(15)
	, DB_SA_I15     =>  DBGSELFADDR0(14)
	, DB_SA_I14     =>  DBGSELFADDR0(13)
	, DB_SA_I13     =>  DBGSELFADDR0(12)
	, DB_SA_I12     =>  DBGSELFADDR0(11)
	, DB_SA_I11     =>  DBGSELFADDR0(10)
	, DB_SA_I10     =>  DBGSELFADDR0(9)
	, DB_SA_I9      =>  DBGSELFADDR0(8)
	, DB_SA_I8      =>  DBGSELFADDR0(7)
	, DB_SA_I7      =>  DBGSELFADDR0(6)
	, DB_SA_I6      =>  DBGSELFADDR0(5)
	, DB_SA_I5      =>  DBGSELFADDR0(4)
	, DB_SA_I4      =>  DBGSELFADDR0(3)
	, DB_SA_I3      =>  DBGSELFADDR0(2)
	, DB_SA_I2      =>  DBGSELFADDR0(1)
	, DB_SA_I1      =>  DBGSELFADDR0(0)

	, DB_SAV_I      =>  DBGSELFADDRV0
	, DEV_E_I       =>  DEVICEEN

	, DFTS_I8       => '0' 
	, DFTS_I7       => '0' 
	, DFTS_I6       => '0' 
	, DFTS_I5       => '0' 
	, DFTS_I4       => '0' 
	, DFTS_I3       => '0' 
	, DFTS_I2       => '0' 
	, DFTS_I1       => '0' 

	, E_DB_I        =>  EDBGRQ0
	, ERR_R_I       =>  ERRENRAM0
	, EVENT_I       =>  EVENTI0

	, GID_I4        =>  GROUPID(3)
	, GID_I3        =>  GROUPID(2)
	, GID_I2        =>  GROUPID(1)
	, GID_I1        =>  GROUPID(0)

	, INIT_P_I      =>  INITPPX0
	, INIT_R_I      =>  INITRAMA0
	, LOC_R_I       =>  LOCZRAMA0
--	, LBK_E_I       =>  LBK_E_I
--	, LBK_MX_I      =>  LBK_MX_I

--	, MODE1_I3      =>  MODE1_I(2)
--	, MODE1_I2      =>  MODE1_I(1)
--	, MODE1_I1      =>  MODE1_I(0)

--	, MODE2_I3      =>  MODE2_I(2)
--	, MODE2_I2      =>  MODE2_I(1)
--	, MODE2_I1      =>  MODE2_I(0)

--	, MODE3_I3      =>  MODE3_I(2)
--	, MODE3_I2      =>  MODE3_I(1)
--	, MODE3_I1      =>  MODE3_I(0)

	, NCPUH_I       =>  nCPUHALT0
	, NET_RS_I      =>  nETMPORESET
	, N_FIQ_I       =>  nFIQ0
	, N_IDE_I       =>  NIDEN0
	, N_IRQ_I       =>  nIRQ0
	, N_PRS_I       =>  nPOTRST
	, N_RS_I        =>  nRESET0
	, N_SPRS_I      =>  nSYSPORESET
	, N_TRS_I       =>  nTRST

	, P_A_I29       =>  PADDRSYS(28)
	, P_A_I28       =>  PADDRSYS(27)
	, P_A_I27       =>  PADDRSYS(26)
	, P_A_I26       =>  PADDRSYS(25)
	, P_A_I25       =>  PADDRSYS(24)
	, P_A_I24       =>  PADDRSYS(23)
	, P_A_I23       =>  PADDRSYS(22)
	, P_A_I22       =>  PADDRSYS(21)
	, P_A_I21       =>  PADDRSYS(20)
	, P_A_I20       =>  PADDRSYS(19)
	, P_A_I19       =>  PADDRSYS(18)
	, P_A_I18       =>  PADDRSYS(17)
	, P_A_I17       =>  PADDRSYS(16)
	, P_A_I16       =>  PADDRSYS(15)
	, P_A_I15       =>  PADDRSYS(14)
	, P_A_I14       =>  PADDRSYS(13)
	, P_A_I13       =>  PADDRSYS(12)
	, P_A_I12       =>  PADDRSYS(11)
	, P_A_I11       =>  PADDRSYS(10)
	, P_A_I10       =>  PADDRSYS(9)
	, P_A_I9        =>  PADDRSYS(8)
	, P_A_I8        =>  PADDRSYS(7)
	, P_A_I7        =>  PADDRSYS(6)
	, P_A_I6        =>  PADDRSYS(5)
	, P_A_I5        =>  PADDRSYS(4)
	, P_A_I4        =>  PADDRSYS(3)
	, P_A_I3        =>  PADDRSYS(2)
	, P_A_I2        =>  PADDRSYS(1)
	, P_A_I1        =>  PADDRSYS(0)

	, P_ECC_I       =>  PARECCENRAM0
	, PLVL_I        =>  PARITYLEVEL
	, P_CK_E_I      =>  PCLKENSYS
	, P_CK_I        =>  PCLKSYS
	, P_E_I         =>  PENABLESYS

	, PPV_BS_I20    =>  PPVBASE0(19)
	, PPV_BS_I19    =>  PPVBASE0(18)
	, PPV_BS_I18    =>  PPVBASE0(17)
	, PPV_BS_I17    =>  PPVBASE0(16)
	, PPV_BS_I16    =>  PPVBASE0(15)
	, PPV_BS_I15    =>  PPVBASE0(14)
	, PPV_BS_I14    =>  PPVBASE0(13)
	, PPV_BS_I13    =>  PPVBASE0(12)
	, PPV_BS_I12    =>  PPVBASE0(11)
	, PPV_BS_I11    =>  PPVBASE0(10)
	, PPV_BS_I10    =>  PPVBASE0(9)
	, PPV_BS_I9     =>  PPVBASE0(8)
	, PPV_BS_I8     =>  PPVBASE0(7)
	, PPV_BS_I7     =>  PPVBASE0(6)
	, PPV_BS_I6     =>  PPVBASE0(5)
	, PPV_BS_I5     =>  PPVBASE0(4)
	, PPV_BS_I4     =>  PPVBASE0(3)
	, PPV_BS_I3     =>  PPVBASE0(2)
	, PPV_BS_I2     =>  PPVBASE0(1)
	, PPV_BS_I1     =>  PPVBASE0(0)

	, PPV_SZ_I5     =>  PPVSIZE0(4)
	, PPV_SZ_I4     =>  PPVSIZE0(3)
	, PPV_SZ_I3     =>  PPVSIZE0(2)
	, PPV_SZ_I2     =>  PPVSIZE0(1)
	, PPV_SZ_I1     =>  PPVSIZE0(0)

	, PPX_BS_I20    =>  PPXBASE0(19)
	, PPX_BS_I19    =>  PPXBASE0(18)
	, PPX_BS_I18    =>  PPXBASE0(17)
	, PPX_BS_I17    =>  PPXBASE0(16)
	, PPX_BS_I16    =>  PPXBASE0(15)
	, PPX_BS_I15    =>  PPXBASE0(14)
	, PPX_BS_I14    =>  PPXBASE0(13)
	, PPX_BS_I13    =>  PPXBASE0(12)
	, PPX_BS_I12    =>  PPXBASE0(11)
	, PPX_BS_I11    =>  PPXBASE0(10)
	, PPX_BS_I10    =>  PPXBASE0(9)
	, PPX_BS_I9     =>  PPXBASE0(8)
	, PPX_BS_I8     =>  PPXBASE0(7)
	, PPX_BS_I7     =>  PPXBASE0(6)
	, PPX_BS_I6     =>  PPXBASE0(5)
	, PPX_BS_I5     =>  PPXBASE0(4)
	, PPX_BS_I4     =>  PPXBASE0(3)
	, PPX_BS_I3     =>  PPXBASE0(2)
	, PPX_BS_I2     =>  PPXBASE0(1)
	, PPX_BS_I1     =>  PPXBASE0(0)

	, PPX_SZ_I5     =>  PPXSIZE0(4)
	, PPX_SZ_I4     =>  PPXSIZE0(3)
	, PPX_SZ_I3     =>  PPXSIZE0(2)
	, PPX_SZ_I2     =>  PPXSIZE0(1)
	, PPX_SZ_I1     =>  PPXSIZE0(0)

	, P_RS_I        =>  PRESETSYSn
	, P_SEL_I       =>  PSELSYS

	, PW_D_I32      =>  PWDATASYS(31)
	, PW_D_I31      =>  PWDATASYS(30)
	, PW_D_I30      =>  PWDATASYS(29)
	, PW_D_I29      =>  PWDATASYS(28)
	, PW_D_I28      =>  PWDATASYS(27)
	, PW_D_I27      =>  PWDATASYS(26)
	, PW_D_I26      =>  PWDATASYS(25)
	, PW_D_I25      =>  PWDATASYS(24)
	, PW_D_I24      =>  PWDATASYS(23)
	, PW_D_I23      =>  PWDATASYS(22)
	, PW_D_I22      =>  PWDATASYS(21)
	, PW_D_I21      =>  PWDATASYS(20)
	, PW_D_I20      =>  PWDATASYS(19)
	, PW_D_I19      =>  PWDATASYS(18)
	, PW_D_I18      =>  PWDATASYS(17)
	, PW_D_I17      =>  PWDATASYS(16)
	, PW_D_I16      =>  PWDATASYS(15)
	, PW_D_I15      =>  PWDATASYS(14)
	, PW_D_I14      =>  PWDATASYS(13)
	, PW_D_I13      =>  PWDATASYS(12)
	, PW_D_I12      =>  PWDATASYS(11)
	, PW_D_I11      =>  PWDATASYS(10)
	, PW_D_I10      =>  PWDATASYS(9)
	, PW_D_I9       =>  PWDATASYS(8)
	, PW_D_I8       =>  PWDATASYS(7)
	, PW_D_I7       =>  PWDATASYS(6)
	, PW_D_I6       =>  PWDATASYS(5)
	, PW_D_I5       =>  PWDATASYS(4)
	, PW_D_I4       =>  PWDATASYS(3)
	, PW_D_I3       =>  PWDATASYS(2)
	, PW_D_I2       =>  PWDATASYS(1)
	, PW_D_I1       =>  PWDATASYS(0)

	, PW_I          =>  PWRITESYS

	, RAMCTL_I8     =>  '0'
	, RAMCTL_I7     =>  '0'
	, RAMCTL_I6     =>  '0'
	, RAMCTL_I5     =>  '0'
	, RAMCTL_I4     =>  '0'
	, RAMCTL_I3     =>  '0'
	, RAMCTL_I2     =>  '0'
	, RAMCTL_I1     =>  '0'

	, R_DM_I64      =>  RDATAM0(63)
	, R_DM_I63      =>  RDATAM0(62)
	, R_DM_I62      =>  RDATAM0(61)
	, R_DM_I61      =>  RDATAM0(60)
	, R_DM_I60      =>  RDATAM0(59)
	, R_DM_I59      =>  RDATAM0(58)
	, R_DM_I58      =>  RDATAM0(57)
	, R_DM_I57      =>  RDATAM0(56)
	, R_DM_I56      =>  RDATAM0(55)
	, R_DM_I55      =>  RDATAM0(54)
	, R_DM_I54      =>  RDATAM0(53)
	, R_DM_I53      =>  RDATAM0(52)
	, R_DM_I52      =>  RDATAM0(51)
	, R_DM_I51      =>  RDATAM0(50)
	, R_DM_I50      =>  RDATAM0(49)
	, R_DM_I49      =>  RDATAM0(48)
	, R_DM_I48      =>  RDATAM0(47)
	, R_DM_I47      =>  RDATAM0(46)
	, R_DM_I46      =>  RDATAM0(45)
	, R_DM_I45      =>  RDATAM0(44)
	, R_DM_I44      =>  RDATAM0(43)
	, R_DM_I43      =>  RDATAM0(42)
	, R_DM_I42      =>  RDATAM0(41)
	, R_DM_I41      =>  RDATAM0(40)
	, R_DM_I40      =>  RDATAM0(39)
	, R_DM_I39      =>  RDATAM0(38)
	, R_DM_I38      =>  RDATAM0(37)
	, R_DM_I37      =>  RDATAM0(36)
	, R_DM_I36      =>  RDATAM0(35)
	, R_DM_I35      =>  RDATAM0(34)
	, R_DM_I34      =>  RDATAM0(33)
	, R_DM_I33      =>  RDATAM0(32)
	, R_DM_I32      =>  RDATAM0(31)
	, R_DM_I31      =>  RDATAM0(30)
	, R_DM_I30      =>  RDATAM0(29)
	, R_DM_I29      =>  RDATAM0(28)
	, R_DM_I28      =>  RDATAM0(27)
	, R_DM_I27      =>  RDATAM0(26)
	, R_DM_I26      =>  RDATAM0(25)
	, R_DM_I25      =>  RDATAM0(24)
	, R_DM_I24      =>  RDATAM0(23)
	, R_DM_I23      =>  RDATAM0(22)
	, R_DM_I22      =>  RDATAM0(21)
	, R_DM_I21      =>  RDATAM0(20)
	, R_DM_I20      =>  RDATAM0(19)
	, R_DM_I19      =>  RDATAM0(18)
	, R_DM_I18      =>  RDATAM0(17)
	, R_DM_I17      =>  RDATAM0(16)
	, R_DM_I16      =>  RDATAM0(15)
	, R_DM_I15      =>  RDATAM0(14)
	, R_DM_I14      =>  RDATAM0(13)
	, R_DM_I13      =>  RDATAM0(12)
	, R_DM_I12      =>  RDATAM0(11)
	, R_DM_I11      =>  RDATAM0(10)
	, R_DM_I10      =>  RDATAM0(9)
	, R_DM_I9       =>  RDATAM0(8)
	, R_DM_I8       =>  RDATAM0(7)
	, R_DM_I7       =>  RDATAM0(6)
	, R_DM_I6       =>  RDATAM0(5)
	, R_DM_I5       =>  RDATAM0(4)
	, R_DM_I4       =>  RDATAM0(3)
	, R_DM_I3       =>  RDATAM0(2)
	, R_DM_I2       =>  RDATAM0(1)
	, R_DM_I1       =>  RDATAM0(0)

	, R_DP_I32      =>  RDATAP0(31)
	, R_DP_I31      =>  RDATAP0(30)
	, R_DP_I30      =>  RDATAP0(29)
	, R_DP_I29      =>  RDATAP0(28)
	, R_DP_I28      =>  RDATAP0(27)
	, R_DP_I27      =>  RDATAP0(26)
	, R_DP_I26      =>  RDATAP0(25)
	, R_DP_I25      =>  RDATAP0(24)
	, R_DP_I24      =>  RDATAP0(23)
	, R_DP_I23      =>  RDATAP0(22)
	, R_DP_I22      =>  RDATAP0(21)
	, R_DP_I21      =>  RDATAP0(20)
	, R_DP_I20      =>  RDATAP0(19)
	, R_DP_I19      =>  RDATAP0(18)
	, R_DP_I18      =>  RDATAP0(17)
	, R_DP_I17      =>  RDATAP0(16)
	, R_DP_I16      =>  RDATAP0(15)
	, R_DP_I15      =>  RDATAP0(14)
	, R_DP_I14      =>  RDATAP0(13)
	, R_DP_I13      =>  RDATAP0(12)
	, R_DP_I12      =>  RDATAP0(11)
	, R_DP_I11      =>  RDATAP0(10)
	, R_DP_I10      =>  RDATAP0(9)
	, R_DP_I9       =>  RDATAP0(8)
	, R_DP_I8       =>  RDATAP0(7)
	, R_DP_I7       =>  RDATAP0(6)
	, R_DP_I6       =>  RDATAP0(5)
	, R_DP_I5       =>  RDATAP0(4)
	, R_DP_I4       =>  RDATAP0(3)
	, R_DP_I3       =>  RDATAP0(2)
	, R_DP_I2       =>  RDATAP0(1)
	, R_DP_I1       =>  RDATAP0(0)

--	, RDY_I3        =>  RDY_I(2)
--	, RDY_I2        =>  RDY_I(1)
--	, RDY_I1        =>  RDY_I(0)

	, R_IDM_I4      =>  RIDM0(3)
	, R_IDM_I3      =>  RIDM0(2)
	, R_IDM_I2      =>  RIDM0(1)
	, R_IDM_I1      =>  RIDM0(0)

	, R_IDP_I4      =>  RIDP0(3)
	, R_IDP_I3      =>  RIDP0(2)
	, R_IDP_I2      =>  RIDP0(1)
	, R_IDP_I1      =>  RIDP0(0)

	, R_LSTM_I      =>  RLASTM0
	, R_LSTP_I      =>  RLASTP0
	, R_RDY_I       =>  RREADYS0

	, R_RSPM_I2     =>  RRESPM0(1)
	, R_RSPM_I1     =>  RRESPM0(0)

	, R_RSPP_I2     =>  RRESPP0(1)
	, R_RSPP_I1     =>  RRESPP0(0)

	, RS_BYP_I      =>  '0'
	, R_VDM_I       =>  RVALIDM0
	, R_VDP_I       =>  RVALIDP0
	, SE_I          =>  '0'
	, SW_CK_I       =>  SWCLKTCK
	, SW_DI_I       =>  SWDITMS
	, T_DI_I        =>  TDI
	, TE_INI_I      =>  TEINIT
	, VINI_I        =>  VINITHI0

	, W_D_I64       =>  WDATAS0(63)
	, W_D_I63       =>  WDATAS0(62)
	, W_D_I62       =>  WDATAS0(61)
	, W_D_I61       =>  WDATAS0(60)
	, W_D_I60       =>  WDATAS0(59)
	, W_D_I59       =>  WDATAS0(58)
	, W_D_I58       =>  WDATAS0(57)
	, W_D_I57       =>  WDATAS0(56)
	, W_D_I56       =>  WDATAS0(55)
	, W_D_I55       =>  WDATAS0(54)
	, W_D_I54       =>  WDATAS0(53)
	, W_D_I53       =>  WDATAS0(52)
	, W_D_I52       =>  WDATAS0(51)
	, W_D_I51       =>  WDATAS0(50)
	, W_D_I50       =>  WDATAS0(49)
	, W_D_I49       =>  WDATAS0(48)
	, W_D_I48       =>  WDATAS0(47)
	, W_D_I47       =>  WDATAS0(46)
	, W_D_I46       =>  WDATAS0(45)
	, W_D_I45       =>  WDATAS0(44)
	, W_D_I44       =>  WDATAS0(43)
	, W_D_I43       =>  WDATAS0(42)
	, W_D_I42       =>  WDATAS0(41)
	, W_D_I41       =>  WDATAS0(40)
	, W_D_I40       =>  WDATAS0(39)
	, W_D_I39       =>  WDATAS0(38)
	, W_D_I38       =>  WDATAS0(37)
	, W_D_I37       =>  WDATAS0(36)
	, W_D_I36       =>  WDATAS0(35)
	, W_D_I35       =>  WDATAS0(34)
	, W_D_I34       =>  WDATAS0(33)
	, W_D_I33       =>  WDATAS0(32)
	, W_D_I32       =>  WDATAS0(31)
	, W_D_I31       =>  WDATAS0(30)
	, W_D_I30       =>  WDATAS0(29)
	, W_D_I29       =>  WDATAS0(28)
	, W_D_I28       =>  WDATAS0(27)
	, W_D_I27       =>  WDATAS0(26)
	, W_D_I26       =>  WDATAS0(25)
	, W_D_I25       =>  WDATAS0(24)
	, W_D_I24       =>  WDATAS0(23)
	, W_D_I23       =>  WDATAS0(22)
	, W_D_I22       =>  WDATAS0(21)
	, W_D_I21       =>  WDATAS0(20)
	, W_D_I20       =>  WDATAS0(19)
	, W_D_I19       =>  WDATAS0(18)
	, W_D_I18       =>  WDATAS0(17)
	, W_D_I17       =>  WDATAS0(16)
	, W_D_I16       =>  WDATAS0(15)
	, W_D_I15       =>  WDATAS0(14)
	, W_D_I14       =>  WDATAS0(13)
	, W_D_I13       =>  WDATAS0(12)
	, W_D_I12       =>  WDATAS0(11)
	, W_D_I11       =>  WDATAS0(10)
	, W_D_I10       =>  WDATAS0(9)
	, W_D_I9        =>  WDATAS0(8)
	, W_D_I8        =>  WDATAS0(7)
	, W_D_I7        =>  WDATAS0(6)
	, W_D_I6        =>  WDATAS0(5)
	, W_D_I5        =>  WDATAS0(4)
	, W_D_I4        =>  WDATAS0(3)
	, W_D_I3        =>  WDATAS0(2)
	, W_D_I2        =>  WDATAS0(1)
	, W_D_I1        =>  WDATAS0(0)

	, W_IDS_I8      =>  WIDS0(7)
	, W_IDS_I7      =>  WIDS0(6)
	, W_IDS_I6      =>  WIDS0(5)
	, W_IDS_I5      =>  WIDS0(4)
	, W_IDS_I4      =>  WIDS0(3)
	, W_IDS_I3      =>  WIDS0(2)
	, W_IDS_I2      =>  WIDS0(1)
	, W_IDS_I1      =>  WIDS0(0)

	, W_LST_I       =>  WLASTS0
	, W_RYM_I       =>  WREADYM0
	, W_RYP_I       =>  WREADYP0

	, W_SBS_I8      =>  WSTRBS0(7)
	, W_SBS_I7      =>  WSTRBS0(6)
	, W_SBS_I6      =>  WSTRBS0(5)
	, W_SBS_I5      =>  WSTRBS0(4)
	, W_SBS_I4      =>  WSTRBS0(3)
	, W_SBS_I3      =>  WSTRBS0(2)
	, W_SBS_I2      =>  WSTRBS0(1)
	, W_SBS_I1      =>  WSTRBS0(0)

	, W_VD_I        =>  WVALIDS0

        -- Outputs
	, AR_AM_O32     =>  ARADDRM0(31)
	, AR_AM_O31     =>  ARADDRM0(30)
	, AR_AM_O30     =>  ARADDRM0(29)
	, AR_AM_O29     =>  ARADDRM0(28)
	, AR_AM_O28     =>  ARADDRM0(27)
	, AR_AM_O27     =>  ARADDRM0(26)
	, AR_AM_O26     =>  ARADDRM0(25)
	, AR_AM_O25     =>  ARADDRM0(24)
	, AR_AM_O24     =>  ARADDRM0(23)
	, AR_AM_O23     =>  ARADDRM0(22)
	, AR_AM_O22     =>  ARADDRM0(21)
	, AR_AM_O21     =>  ARADDRM0(20)
	, AR_AM_O20     =>  ARADDRM0(19)
	, AR_AM_O19     =>  ARADDRM0(18)
	, AR_AM_O18     =>  ARADDRM0(17)
	, AR_AM_O17     =>  ARADDRM0(16)
	, AR_AM_O16     =>  ARADDRM0(15)
	, AR_AM_O15     =>  ARADDRM0(14)
	, AR_AM_O14     =>  ARADDRM0(13)
	, AR_AM_O13     =>  ARADDRM0(12)
	, AR_AM_O12     =>  ARADDRM0(11)
	, AR_AM_O11     =>  ARADDRM0(10)
	, AR_AM_O10     =>  ARADDRM0(9)
	, AR_AM_O9      =>  ARADDRM0(8)
	, AR_AM_O8      =>  ARADDRM0(7)
	, AR_AM_O7      =>  ARADDRM0(6)
	, AR_AM_O6      =>  ARADDRM0(5)
	, AR_AM_O5      =>  ARADDRM0(4)
	, AR_AM_O4      =>  ARADDRM0(3)
	, AR_AM_O3      =>  ARADDRM0(2)
	, AR_AM_O2      =>  ARADDRM0(1)
	, AR_AM_O1      =>  ARADDRM0(0)

	, AR_AP_O32     =>  ARADDRP0(31)
	, AR_AP_O31     =>  ARADDRP0(30)
	, AR_AP_O30     =>  ARADDRP0(29)
	, AR_AP_O29     =>  ARADDRP0(28)
	, AR_AP_O28     =>  ARADDRP0(27)
	, AR_AP_O27     =>  ARADDRP0(26)
	, AR_AP_O26     =>  ARADDRP0(25)
	, AR_AP_O25     =>  ARADDRP0(24)
	, AR_AP_O24     =>  ARADDRP0(23)
	, AR_AP_O23     =>  ARADDRP0(22)
	, AR_AP_O22     =>  ARADDRP0(21)
	, AR_AP_O21     =>  ARADDRP0(20)
	, AR_AP_O20     =>  ARADDRP0(19)
	, AR_AP_O19     =>  ARADDRP0(18)
	, AR_AP_O18     =>  ARADDRP0(17)
	, AR_AP_O17     =>  ARADDRP0(16)
	, AR_AP_O16     =>  ARADDRP0(15)
	, AR_AP_O15     =>  ARADDRP0(14)
	, AR_AP_O14     =>  ARADDRP0(13)
	, AR_AP_O13     =>  ARADDRP0(12)
	, AR_AP_O12     =>  ARADDRP0(11)
	, AR_AP_O11     =>  ARADDRP0(10)
	, AR_AP_O10     =>  ARADDRP0(9)
	, AR_AP_O9      =>  ARADDRP0(8)
	, AR_AP_O8      =>  ARADDRP0(7)
	, AR_AP_O7      =>  ARADDRP0(6)
	, AR_AP_O6      =>  ARADDRP0(5)
	, AR_AP_O5      =>  ARADDRP0(4)
	, AR_AP_O4      =>  ARADDRP0(3)
	, AR_AP_O3      =>  ARADDRP0(2)
	, AR_AP_O2      =>  ARADDRP0(1)
	, AR_AP_O1      =>  ARADDRP0(0)

	, AR_BUM_O2     =>  ARBURSTM0(1)
	, AR_BUM_O1     =>  ARBURSTM0(0)

	, AR_BUP_O2     =>  ARBURSTP0(1)
	, AR_BUP_O1     =>  ARBURSTP0(0)

	, AR_CHM_O4     =>  ARCACHEM0(3)
	, AR_CHM_O3     =>  ARCACHEM0(2)
	, AR_CHM_O2     =>  ARCACHEM0(1)
	, AR_CHM_O1     =>  ARCACHEM0(0)

	, AR_CHP_O4     =>  ARCACHEP0(3)
	, AR_CHP_O3     =>  ARCACHEP0(2)
	, AR_CHP_O2     =>  ARCACHEP0(1)
	, AR_CHP_O1     =>  ARCACHEP0(0)

	, AR_IDM_O4     =>  ARIDM0(3)
	, AR_IDM_O3     =>  ARIDM0(2)
	, AR_IDM_O2     =>  ARIDM0(1)
	, AR_IDM_O1     =>  ARIDM0(0)

	, AR_IDP_O4     =>  ARIDP0(3)
	, AR_IDP_O3     =>  ARIDP0(2)
	, AR_IDP_O2     =>  ARIDP0(1)
	, AR_IDP_O1     =>  ARIDP0(0)

	, AR_INM_O4     =>  ARINNERM0(3)
	, AR_INM_O3     =>  ARINNERM0(2)
	, AR_INM_O2     =>  ARINNERM0(1)
	, AR_INM_O1     =>  ARINNERM0(0)

	, AR_LEM_O4     =>  ARLENM0(3)
	, AR_LEM_O3     =>  ARLENM0(2)
	, AR_LEM_O2     =>  ARLENM0(1)
	, AR_LEM_O1     =>  ARLENM0(0)

	, AR_LEP_O4     =>  ARLENP0(3)
	, AR_LEP_O3     =>  ARLENP0(2)
	, AR_LEP_O2     =>  ARLENP0(1)
	, AR_LEP_O1     =>  ARLENP0(0)

	, AR_LKM_O2     =>  ARLOCKM0(1)
	, AR_LKM_O1     =>  ARLOCKM0(0)

	, AR_LKP_O2     =>  ARLOCKP0(1)
	, AR_LKP_O1     =>  ARLOCKP0(0)

	, AR_PRM_O3     =>  ARPROTM0(2)
	, AR_PRM_O2     =>  ARPROTM0(1)
	, AR_PRM_O1     =>  ARPROTM0(0)

	, AR_PRP_O3     =>  ARPROTP0(2)
	, AR_PRP_O2     =>  ARPROTP0(1)
	, AR_PRP_O1     =>  ARPROTP0(0)

	, AR_RDY_O      =>  ARREADYS0
	, AR_SHM_O      =>  ARSHAREM0

	, AR_SZM_O3     =>  ARSIZEM0(2)
	, AR_SZM_O2     =>  ARSIZEM0(1)
	, AR_SZM_O1     =>  ARSIZEM0(0)

	, AR_SZP_O3     =>  ARSIZEP0(2)
	, AR_SZP_O2     =>  ARSIZEP0(1)
	, AR_SZP_O1     =>  ARSIZEP0(0)

	, AR_VDM_O      =>  ARVALIDM0
	, AR_VDP_O      =>  ARVALIDP0

	, AW_AM_O32     =>  AWADDRM0(31)
	, AW_AM_O31     =>  AWADDRM0(30)
	, AW_AM_O30     =>  AWADDRM0(29)
	, AW_AM_O29     =>  AWADDRM0(28)
	, AW_AM_O28     =>  AWADDRM0(27)
	, AW_AM_O27     =>  AWADDRM0(26)
	, AW_AM_O26     =>  AWADDRM0(25)
	, AW_AM_O25     =>  AWADDRM0(24)
	, AW_AM_O24     =>  AWADDRM0(23)
	, AW_AM_O23     =>  AWADDRM0(22)
	, AW_AM_O22     =>  AWADDRM0(21)
	, AW_AM_O21     =>  AWADDRM0(20)
	, AW_AM_O20     =>  AWADDRM0(19)
	, AW_AM_O19     =>  AWADDRM0(18)
	, AW_AM_O18     =>  AWADDRM0(17)
	, AW_AM_O17     =>  AWADDRM0(16)
	, AW_AM_O16     =>  AWADDRM0(15)
	, AW_AM_O15     =>  AWADDRM0(14)
	, AW_AM_O14     =>  AWADDRM0(13)
	, AW_AM_O13     =>  AWADDRM0(12)
	, AW_AM_O12     =>  AWADDRM0(11)
	, AW_AM_O11     =>  AWADDRM0(10)
	, AW_AM_O10     =>  AWADDRM0(9)
	, AW_AM_O9      =>  AWADDRM0(8)
	, AW_AM_O8      =>  AWADDRM0(7)
	, AW_AM_O7      =>  AWADDRM0(6)
	, AW_AM_O6      =>  AWADDRM0(5)
	, AW_AM_O5      =>  AWADDRM0(4)
	, AW_AM_O4      =>  AWADDRM0(3)
	, AW_AM_O3      =>  AWADDRM0(2)
	, AW_AM_O2      =>  AWADDRM0(1)
	, AW_AM_O1      =>  AWADDRM0(0)

	, AW_AP_O32     =>  AWADDRP0(31)
	, AW_AP_O31     =>  AWADDRP0(30)
	, AW_AP_O30     =>  AWADDRP0(29)
	, AW_AP_O29     =>  AWADDRP0(28)
	, AW_AP_O28     =>  AWADDRP0(27)
	, AW_AP_O27     =>  AWADDRP0(26)
	, AW_AP_O26     =>  AWADDRP0(25)
	, AW_AP_O25     =>  AWADDRP0(24)
	, AW_AP_O24     =>  AWADDRP0(23)
	, AW_AP_O23     =>  AWADDRP0(22)
	, AW_AP_O22     =>  AWADDRP0(21)
	, AW_AP_O21     =>  AWADDRP0(20)
	, AW_AP_O20     =>  AWADDRP0(19)
	, AW_AP_O19     =>  AWADDRP0(18)
	, AW_AP_O18     =>  AWADDRP0(17)
	, AW_AP_O17     =>  AWADDRP0(16)
	, AW_AP_O16     =>  AWADDRP0(15)
	, AW_AP_O15     =>  AWADDRP0(14)
	, AW_AP_O14     =>  AWADDRP0(13)
	, AW_AP_O13     =>  AWADDRP0(12)
	, AW_AP_O12     =>  AWADDRP0(11)
	, AW_AP_O11     =>  AWADDRP0(10)
	, AW_AP_O10     =>  AWADDRP0(9)
	, AW_AP_O9      =>  AWADDRP0(8)
	, AW_AP_O8      =>  AWADDRP0(7)
	, AW_AP_O7      =>  AWADDRP0(6)
	, AW_AP_O6      =>  AWADDRP0(5)
	, AW_AP_O5      =>  AWADDRP0(4)
	, AW_AP_O4      =>  AWADDRP0(3)
	, AW_AP_O3      =>  AWADDRP0(2)
	, AW_AP_O2      =>  AWADDRP0(1)
	, AW_AP_O1      =>  AWADDRP0(0)

	, AW_BUM_O2     =>  AWBURSTM0(1)
	, AW_BUM_O1     =>  AWBURSTM0(0)

	, AW_BUP_O2     =>  AWBURSTP0(1)
	, AW_BUP_O1     =>  AWBURSTP0(0)

	, AW_CHM_O4     =>  AWCACHEM0(3)
	, AW_CHM_O3     =>  AWCACHEM0(2)
	, AW_CHM_O2     =>  AWCACHEM0(1)
	, AW_CHM_O1     =>  AWCACHEM0(0)

	, AW_CHP_O4     =>  AWCACHEP0(3)
	, AW_CHP_O3     =>  AWCACHEP0(2)
	, AW_CHP_O2     =>  AWCACHEP0(1)
	, AW_CHP_O1     =>  AWCACHEP0(0)

	, AW_IDM_O4     =>  AWIDM0(3)
	, AW_IDM_O3     =>  AWIDM0(2)
	, AW_IDM_O2     =>  AWIDM0(1)
	, AW_IDM_O1     =>  AWIDM0(0)

	, AW_IDP_O4     =>  AWIDP0(3)
	, AW_IDP_O3     =>  AWIDP0(2)
	, AW_IDP_O2     =>  AWIDP0(1)
	, AW_IDP_O1     =>  AWIDP0(0)

	, AW_INM_O4     =>  AWINNERM0(3)
	, AW_INM_O3     =>  AWINNERM0(2)
	, AW_INM_O2     =>  AWINNERM0(1)
	, AW_INM_O1     =>  AWINNERM0(0)

	, AW_LEM_O4     =>  AWLENM0(3)
	, AW_LEM_O3     =>  AWLENM0(2)
	, AW_LEM_O2     =>  AWLENM0(1)
	, AW_LEM_O1     =>  AWLENM0(0)

	, AW_LEP_O4     =>  AWLENP0(3)
	, AW_LEP_O3     =>  AWLENP0(2)
	, AW_LEP_O2     =>  AWLENP0(1)
	, AW_LEP_O1     =>  AWLENP0(0)

	, AW_LKM_O2     =>  AWLOCKM0(1)
	, AW_LKM_O1     =>  AWLOCKM0(0)

	, AW_LKP_O2     =>  AWLOCKP0(1)
	, AW_LKP_O1     =>  AWLOCKP0(0)

	, AW_PRM_O3     =>  AWPROTM0(2)
	, AW_PRM_O2     =>  AWPROTM0(1)
	, AW_PRM_O1     =>  AWPROTM0(0)

	, AW_PRP_O3     =>  AWPROTP0(2)
	, AW_PRP_O2     =>  AWPROTP0(1)
	, AW_PRP_O1     =>  AWPROTP0(0)

	, AW_RDY_O      =>  AWREADYS0
	, AW_SHM_O      =>  AWSHAREM0

	, AW_SZM_O3     =>  AWSIZEM0(2)
	, AW_SZM_O2     =>  AWSIZEM0(1)
	, AW_SZM_O1     =>  AWSIZEM0(0)

	, AW_SZP_O3     =>  AWSIZEP0(2)
	, AW_SZP_O2     =>  AWSIZEP0(1)
	, AW_SZP_O1     =>  AWSIZEP0(0)

	, AW_VDM_O      =>  AWVALIDM0
	, AW_VDP_O      =>  AWVALIDP0

	, B_IDS_O8      =>  BIDS0(7)
	, B_IDS_O7      =>  BIDS0(6)
	, B_IDS_O6      =>  BIDS0(5)
	, B_IDS_O5      =>  BIDS0(4)
	, B_IDS_O4      =>  BIDS0(3)
	, B_IDS_O3      =>  BIDS0(2)
	, B_IDS_O2      =>  BIDS0(1)
	, B_IDS_O1      =>  BIDS0(0)

	, B_RDYM_O      =>  BREADYM0
	, B_RDYP_O      =>  BREADYP0

	, B_RSP_O2      =>  BRESPS0(1)
	, B_RSP_O1      =>  BRESPS0(0)

	, B_VD_O        =>  BVALIDS0

	, CDB_PW_O      =>  CDBGPWRUPREQ
	, CDB_RS_O      =>  CDBGRSTREQ
	, COM_RX_O      =>  COMMRX0
	, COM_TX_O      =>  COMMTX0
	, CS_PW_O       =>  CSYSPWRUPREQ
	, DB_ACK_O      =>  DBGACK0
	, DB_NPD_O      =>  DBGNOPWRDWN
	, DB_RS_O       =>  DBGRSTREQ0

	, DFTS_O8       =>  open
	, DFTS_O7       =>  open
	, DFTS_O6       =>  open
	, DFTS_O5       =>  open
	, DFTS_O4       =>  open
	, DFTS_O3       =>  open
	, DFTS_O2       =>  open
	, DFTS_O1       =>  open

	, ET_ASC_O8     =>  ETMASICCTL0(7)
	, ET_ASC_O7     =>  ETMASICCTL0(6)
	, ET_ASC_O6     =>  ETMASICCTL0(5)
	, ET_ASC_O5     =>  ETMASICCTL0(4)
	, ET_ASC_O4     =>  ETMASICCTL0(3)
	, ET_ASC_O3     =>  ETMASICCTL0(2)
	, ET_ASC_O2     =>  ETMASICCTL0(1)
	, ET_ASC_O1     =>  ETMASICCTL0(0)

	, ET_E_O        =>  ETMEN0

	, ET_EXT_O2     =>  ETMEXTOUT0(1)
	, ET_EXT_O1     =>  ETMEXTOUT0(0)

	, EVENT_O       =>  EVENTO0
	, FP_DZC_O      =>  FPDZC0
	, FP_IDC_O      =>  FPIDC0
	, FP_IOC_O      =>  FPIOC0
	, FP_IXC_O      =>  FPIXC0
	, FP_OFC_O      =>  FPOFC0
	, FP_UFC_O      =>  FPUFC0
	, JTAG_O        =>  JTAGNSW


	, N_CKST_O      =>  nCLKSTOPPED0
	, N_PMU_O       =>  nPMUIRQ0
	, N_TDO_O       =>  nTDOEN
	, N_VFIQ_O      =>  nVALFIQ0
	, N_VIRQ_O      =>  nVALIRQ0
	, N_VRST_O      =>  nVALRESET0
	, N_EPST_O      =>  nWFEPIPESTOPPED0
	, N_IPST_O      =>  nWFIPIPESTOPPED0

	, P_RD_O32      =>  PRDATASYS(31)
	, P_RD_O31      =>  PRDATASYS(30)
	, P_RD_O30      =>  PRDATASYS(29)
	, P_RD_O29      =>  PRDATASYS(28)
	, P_RD_O28      =>  PRDATASYS(27)
	, P_RD_O27      =>  PRDATASYS(26)
	, P_RD_O26      =>  PRDATASYS(25)
	, P_RD_O25      =>  PRDATASYS(24)
	, P_RD_O24      =>  PRDATASYS(23)
	, P_RD_O23      =>  PRDATASYS(22)
	, P_RD_O22      =>  PRDATASYS(21)
	, P_RD_O21      =>  PRDATASYS(20)
	, P_RD_O20      =>  PRDATASYS(19)
	, P_RD_O19      =>  PRDATASYS(18)
	, P_RD_O18      =>  PRDATASYS(17)
	, P_RD_O17      =>  PRDATASYS(16)
	, P_RD_O16      =>  PRDATASYS(15)
	, P_RD_O15      =>  PRDATASYS(14)
	, P_RD_O14      =>  PRDATASYS(13)
	, P_RD_O13      =>  PRDATASYS(12)
	, P_RD_O12      =>  PRDATASYS(11)
	, P_RD_O11      =>  PRDATASYS(10)
	, P_RD_O10      =>  PRDATASYS(9)
	, P_RD_O9       =>  PRDATASYS(8)
	, P_RD_O8       =>  PRDATASYS(7)
	, P_RD_O7       =>  PRDATASYS(6)
	, P_RD_O6       =>  PRDATASYS(5)
	, P_RD_O5       =>  PRDATASYS(4)
	, P_RD_O4       =>  PRDATASYS(3)
	, P_RD_O3       =>  PRDATASYS(2)
	, P_RD_O2       =>  PRDATASYS(1)
	, P_RD_O1       =>  PRDATASYS(0)

	, P_RDY_O       =>  PREADYSYS
	, P_VER_O       =>  PSLVERRSYS

	, RD_O64        =>  RDATAS0(63)
	, RD_O63        =>  RDATAS0(62)
	, RD_O62        =>  RDATAS0(61)
	, RD_O61        =>  RDATAS0(60)
	, RD_O60        =>  RDATAS0(59)
	, RD_O59        =>  RDATAS0(58)
	, RD_O58        =>  RDATAS0(57)
	, RD_O57        =>  RDATAS0(56)
	, RD_O56        =>  RDATAS0(55)
	, RD_O55        =>  RDATAS0(54)
	, RD_O54        =>  RDATAS0(53)
	, RD_O53        =>  RDATAS0(52)
	, RD_O52        =>  RDATAS0(51)
	, RD_O51        =>  RDATAS0(50)
	, RD_O50        =>  RDATAS0(49)
	, RD_O49        =>  RDATAS0(48)
	, RD_O48        =>  RDATAS0(47)
	, RD_O47        =>  RDATAS0(46)
	, RD_O46        =>  RDATAS0(45)
	, RD_O45        =>  RDATAS0(44)
	, RD_O44        =>  RDATAS0(43)
	, RD_O43        =>  RDATAS0(42)
	, RD_O42        =>  RDATAS0(41)
	, RD_O41        =>  RDATAS0(40)
	, RD_O40        =>  RDATAS0(39)
	, RD_O39        =>  RDATAS0(38)
	, RD_O38        =>  RDATAS0(37)
	, RD_O37        =>  RDATAS0(36)
	, RD_O36        =>  RDATAS0(35)
	, RD_O35        =>  RDATAS0(34)
	, RD_O34        =>  RDATAS0(33)
	, RD_O33        =>  RDATAS0(32)
	, RD_O32        =>  RDATAS0(31)
	, RD_O31        =>  RDATAS0(30)
	, RD_O30        =>  RDATAS0(29)
	, RD_O29        =>  RDATAS0(28)
	, RD_O28        =>  RDATAS0(27)
	, RD_O27        =>  RDATAS0(26)
	, RD_O26        =>  RDATAS0(25)
	, RD_O25        =>  RDATAS0(24)
	, RD_O24        =>  RDATAS0(23)
	, RD_O23        =>  RDATAS0(22)
	, RD_O22        =>  RDATAS0(21)
	, RD_O21        =>  RDATAS0(20)
	, RD_O20        =>  RDATAS0(19)
	, RD_O19        =>  RDATAS0(18)
	, RD_O18        =>  RDATAS0(17)
	, RD_O17        =>  RDATAS0(16)
	, RD_O16        =>  RDATAS0(15)
	, RD_O15        =>  RDATAS0(14)
	, RD_O14        =>  RDATAS0(13)
	, RD_O13        =>  RDATAS0(12)
	, RD_O12        =>  RDATAS0(11)
	, RD_O11        =>  RDATAS0(10)
	, RD_O10        =>  RDATAS0(9)
	, RD_O9         =>  RDATAS0(8)
	, RD_O8         =>  RDATAS0(7)
	, RD_O7         =>  RDATAS0(6)
	, RD_O6         =>  RDATAS0(5)
	, RD_O5         =>  RDATAS0(4)
	, RD_O4         =>  RDATAS0(3)
	, RD_O3         =>  RDATAS0(2)
	, RD_O2         =>  RDATAS0(1)
	, RD_O1         =>  RDATAS0(0)



	, R_IDS_O8      =>  RIDS0(7)
	, R_IDS_O7      =>  RIDS0(6)
	, R_IDS_O6      =>  RIDS0(5)
	, R_IDS_O5      =>  RIDS0(4)
	, R_IDS_O4      =>  RIDS0(3)
	, R_IDS_O3      =>  RIDS0(2)
	, R_IDS_O2      =>  RIDS0(1)
	, R_IDS_O1      =>  RIDS0(0)

	, R_LST_O       =>  RLASTS0
	, R_RDYM_O      =>  RREADYM0
	, R_RDYP_O      =>  RREADYP0

	, R_RSP_O2      =>  RRESPS0(1)
	, R_RSP_O1      =>  RRESPS0(0)

	, R_VD_O        =>  RVALIDS0

	, SWDO_O        =>  SWDO
	, SWDO_E_O      =>  SWDOEN
	, TDO_O         =>  TDO
	, T_CK_O        =>  TRACECLK
	, T_CTL_O       =>  TRACECTL

	, T_DATA_O32    =>  TRACEDATA(31)
	, T_DATA_O31    =>  TRACEDATA(30)
	, T_DATA_O30    =>  TRACEDATA(29)
	, T_DATA_O29    =>  TRACEDATA(28)
	, T_DATA_O28    =>  TRACEDATA(27)
	, T_DATA_O27    =>  TRACEDATA(26)
	, T_DATA_O26    =>  TRACEDATA(25)
	, T_DATA_O25    =>  TRACEDATA(24)
	, T_DATA_O24    =>  TRACEDATA(23)
	, T_DATA_O23    =>  TRACEDATA(22)
	, T_DATA_O22    =>  TRACEDATA(21)
	, T_DATA_O21    =>  TRACEDATA(20)
	, T_DATA_O20    =>  TRACEDATA(19)
	, T_DATA_O19    =>  TRACEDATA(18)
	, T_DATA_O18    =>  TRACEDATA(17)
	, T_DATA_O17    =>  TRACEDATA(16)
	, T_DATA_O16    =>  TRACEDATA(15)
	, T_DATA_O15    =>  TRACEDATA(14)
	, T_DATA_O14    =>  TRACEDATA(13)
	, T_DATA_O13    =>  TRACEDATA(12)
	, T_DATA_O12    =>  TRACEDATA(11)
	, T_DATA_O11    =>  TRACEDATA(10)
	, T_DATA_O10    =>  TRACEDATA(9)
	, T_DATA_O9     =>  TRACEDATA(8)
	, T_DATA_O8     =>  TRACEDATA(7)
	, T_DATA_O7     =>  TRACEDATA(6)
	, T_DATA_O6     =>  TRACEDATA(5)
	, T_DATA_O5     =>  TRACEDATA(4)
	, T_DATA_O4     =>  TRACEDATA(3)
	, T_DATA_O3     =>  TRACEDATA(2)
	, T_DATA_O2     =>  TRACEDATA(1)
	, T_DATA_O1     =>  TRACEDATA(0)


	, W_DM_O64      =>  WDATAM0(63)
	, W_DM_O63      =>  WDATAM0(62)
	, W_DM_O62      =>  WDATAM0(61)
	, W_DM_O61      =>  WDATAM0(60)
	, W_DM_O60      =>  WDATAM0(59)
	, W_DM_O59      =>  WDATAM0(58)
	, W_DM_O58      =>  WDATAM0(57)
	, W_DM_O57      =>  WDATAM0(56)
	, W_DM_O56      =>  WDATAM0(55)
	, W_DM_O55      =>  WDATAM0(54)
	, W_DM_O54      =>  WDATAM0(53)
	, W_DM_O53      =>  WDATAM0(52)
	, W_DM_O52      =>  WDATAM0(51)
	, W_DM_O51      =>  WDATAM0(50)
	, W_DM_O50      =>  WDATAM0(49)
	, W_DM_O49      =>  WDATAM0(48)
	, W_DM_O48      =>  WDATAM0(47)
	, W_DM_O47      =>  WDATAM0(46)
	, W_DM_O46      =>  WDATAM0(45)
	, W_DM_O45      =>  WDATAM0(44)
	, W_DM_O44      =>  WDATAM0(43)
	, W_DM_O43      =>  WDATAM0(42)
	, W_DM_O42      =>  WDATAM0(41)
	, W_DM_O41      =>  WDATAM0(40)
	, W_DM_O40      =>  WDATAM0(39)
	, W_DM_O39      =>  WDATAM0(38)
	, W_DM_O38      =>  WDATAM0(37)
	, W_DM_O37      =>  WDATAM0(36)
	, W_DM_O36      =>  WDATAM0(35)
	, W_DM_O35      =>  WDATAM0(34)
	, W_DM_O34      =>  WDATAM0(33)
	, W_DM_O33      =>  WDATAM0(32)
	, W_DM_O32      =>  WDATAM0(31)
	, W_DM_O31      =>  WDATAM0(30)
	, W_DM_O30      =>  WDATAM0(29)
	, W_DM_O29      =>  WDATAM0(28)
	, W_DM_O28      =>  WDATAM0(27)
	, W_DM_O27      =>  WDATAM0(26)
	, W_DM_O26      =>  WDATAM0(25)
	, W_DM_O25      =>  WDATAM0(24)
	, W_DM_O24      =>  WDATAM0(23)
	, W_DM_O23      =>  WDATAM0(22)
	, W_DM_O22      =>  WDATAM0(21)
	, W_DM_O21      =>  WDATAM0(20)
	, W_DM_O20      =>  WDATAM0(19)
	, W_DM_O19      =>  WDATAM0(18)
	, W_DM_O18      =>  WDATAM0(17)
	, W_DM_O17      =>  WDATAM0(16)
	, W_DM_O16      =>  WDATAM0(15)
	, W_DM_O15      =>  WDATAM0(14)
	, W_DM_O14      =>  WDATAM0(13)
	, W_DM_O13      =>  WDATAM0(12)
	, W_DM_O12      =>  WDATAM0(11)
	, W_DM_O11      =>  WDATAM0(10)
	, W_DM_O10      =>  WDATAM0(9)
	, W_DM_O9       =>  WDATAM0(8)
	, W_DM_O8       =>  WDATAM0(7)
	, W_DM_O7       =>  WDATAM0(6)
	, W_DM_O6       =>  WDATAM0(5)
	, W_DM_O5       =>  WDATAM0(4)
	, W_DM_O4       =>  WDATAM0(3)
	, W_DM_O3       =>  WDATAM0(2)
	, W_DM_O2       =>  WDATAM0(1)
	, W_DM_O1       =>  WDATAM0(0)

	, W_DP_O32      =>  WDATAP0(31)
	, W_DP_O31      =>  WDATAP0(30)
	, W_DP_O30      =>  WDATAP0(29)
	, W_DP_O29      =>  WDATAP0(28)
	, W_DP_O28      =>  WDATAP0(27)
	, W_DP_O27      =>  WDATAP0(26)
	, W_DP_O26      =>  WDATAP0(25)
	, W_DP_O25      =>  WDATAP0(24)
	, W_DP_O24      =>  WDATAP0(23)
	, W_DP_O23      =>  WDATAP0(22)
	, W_DP_O22      =>  WDATAP0(21)
	, W_DP_O21      =>  WDATAP0(20)
	, W_DP_O20      =>  WDATAP0(19)
	, W_DP_O19      =>  WDATAP0(18)
	, W_DP_O18      =>  WDATAP0(17)
	, W_DP_O17      =>  WDATAP0(16)
	, W_DP_O16      =>  WDATAP0(15)
	, W_DP_O15      =>  WDATAP0(14)
	, W_DP_O14      =>  WDATAP0(13)
	, W_DP_O13      =>  WDATAP0(12)
	, W_DP_O12      =>  WDATAP0(11)
	, W_DP_O11      =>  WDATAP0(10)
	, W_DP_O10      =>  WDATAP0(9)
	, W_DP_O9       =>  WDATAP0(8)
	, W_DP_O8       =>  WDATAP0(7)
	, W_DP_O7       =>  WDATAP0(6)
	, W_DP_O6       =>  WDATAP0(5)
	, W_DP_O5       =>  WDATAP0(4)
	, W_DP_O4       =>  WDATAP0(3)
	, W_DP_O3       =>  WDATAP0(2)
	, W_DP_O2       =>  WDATAP0(1)
	, W_DP_O1       =>  WDATAP0(0)

	, W_IDM_O4      =>  WIDM0(3)
	, W_IDM_O3      =>  WIDM0(2)
	, W_IDM_O2      =>  WIDM0(1)
	, W_IDM_O1      =>  WIDM0(0)

	, W_IDP_O4      =>  WIDP0(3)
	, W_IDP_O3      =>  WIDP0(2)
	, W_IDP_O2      =>  WIDP0(1)
	, W_IDP_O1      =>  WIDP0(0)

	, W_LSTM_O      =>  WLASTM0
	, W_LSTP_O      =>  WLASTP0
	, W_RDY_O       =>  WREADYS0

	, W_SBM_O8      =>  WSTRBM0(7)
	, W_SBM_O7      =>  WSTRBM0(6)
	, W_SBM_O6      =>  WSTRBM0(5)
	, W_SBM_O5      =>  WSTRBM0(4)
	, W_SBM_O4      =>  WSTRBM0(3)
	, W_SBM_O3      =>  WSTRBM0(2)
	, W_SBM_O2      =>  WSTRBM0(1)
	, W_SBM_O1      =>  WSTRBM0(0)

	, W_SBP_O4      =>  WSTRBP0(3)
	, W_SBP_O3      =>  WSTRBP0(2)
	, W_SBP_O2      =>  WSTRBP0(1)
	, W_SBP_O1      =>  WSTRBP0(0)

	, W_VDM_O       =>  WVALIDM0
	, W_VDP_O       =>  WVALIDP0
);
end NX_RTL;
-- =================================================================================================
--   NX_RB definition                                                                   2020/04/08
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_RB is
generic (
    -- input : EI to FO
    inputClk      : bit_vector( 1 downto 0) := B"00"; -- 00 = CK1, 01 = CK2, 10 = CK3 and 11 = CK4
    inputBypass   : bit_vector(23 downto 0) := B"000000000000000000000000"; -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    inputContext  : string := ""; -- input context initialization
    -- output : FI to EO
    outputClk     : bit_vector( 1 downto 0) := B"00"; -- 00 = CK1, 01 = CK2, 10 = CK3 and 11 = CK4
    outputBypass  : bit_vector(23 downto 0) := B"000000000000000000000000";  -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    outputContext : string := "" -- output context initialization
);
port (
    CK1   : in  std_logic;
    CK2   : in  std_logic;
    CK3   : in  std_logic;
    CK4   : in  std_logic;
    EI1   : in  std_logic;
    EI2   : in  std_logic;
    EI3   : in  std_logic;
    EI4   : in  std_logic;
    EI5   : in  std_logic;
    EI6   : in  std_logic;
    EI7   : in  std_logic;
    EI8   : in  std_logic;
    EI9   : in  std_logic;
    EI10  : in  std_logic;
    EI11  : in  std_logic;
    EI12  : in  std_logic;
    EI13  : in  std_logic;
    EI14  : in  std_logic;
    EI15  : in  std_logic;
    EI16  : in  std_logic;
    EI17  : in  std_logic;
    EI18  : in  std_logic;
    EI19  : in  std_logic;
    EI20  : in  std_logic;
    EI21  : in  std_logic;
    EI22  : in  std_logic;
    EI23  : in  std_logic;
    EI24  : in  std_logic;
    EI25  : in  std_logic;
    EI26  : in  std_logic;
    EI27  : in  std_logic;
    EI28  : in  std_logic;
    EI29  : in  std_logic;
    EI30  : in  std_logic;
    EI31  : in  std_logic;
    EI32  : in  std_logic;
    EI33  : in  std_logic;
    EI34  : in  std_logic;
    EI35  : in  std_logic;
    EI36  : in  std_logic;
    EI37  : in  std_logic;
    EI38  : in  std_logic;
    EI39  : in  std_logic;
    EI40  : in  std_logic;
    EI41  : in  std_logic;
    EI42  : in  std_logic;
    EI43  : in  std_logic;
    EI44  : in  std_logic;
    EI45  : in  std_logic;
    EI46  : in  std_logic;
    EI47  : in  std_logic;
    EI48  : in  std_logic;
    EI49  : in  std_logic;
    EI50  : in  std_logic;
    EI51  : in  std_logic;
    EI52  : in  std_logic;
    EI53  : in  std_logic;
    EI54  : in  std_logic;
    EI55  : in  std_logic;
    EI56  : in  std_logic;
    EI57  : in  std_logic;
    EI58  : in  std_logic;
    EI59  : in  std_logic;
    EI60  : in  std_logic;
    EI61  : in  std_logic;
    EI62  : in  std_logic;
    EI63  : in  std_logic;
    EI64  : in  std_logic;
    EI65  : in  std_logic;
    EI66  : in  std_logic;
    EI67  : in  std_logic;
    EI68  : in  std_logic;
    EI69  : in  std_logic;
    EI70  : in  std_logic;
    EI71  : in  std_logic;
    EI72  : in  std_logic;
    EI73  : in  std_logic;
    EI74  : in  std_logic;
    EI75  : in  std_logic;
    EI76  : in  std_logic;
    EI77  : in  std_logic;
    EI78  : in  std_logic;
    EI79  : in  std_logic;
    EI80  : in  std_logic;
    EI81  : in  std_logic;
    EI82  : in  std_logic;
    EI83  : in  std_logic;
    EI84  : in  std_logic;
    EI85  : in  std_logic;
    EI86  : in  std_logic;
    EI87  : in  std_logic;
    EI88  : in  std_logic;
    EI89  : in  std_logic;
    EI90  : in  std_logic;
    EI91  : in  std_logic;
    EI92  : in  std_logic;
    EI93  : in  std_logic;
    EI94  : in  std_logic;
    EI95  : in  std_logic;
    EI96  : in  std_logic;
    EI97  : in  std_logic;
    EI98  : in  std_logic;
    EI99  : in  std_logic;
    EI100 : in  std_logic;
    EI101 : in  std_logic;
    EI102 : in  std_logic;
    EI103 : in  std_logic;
    EI104 : in  std_logic;
    EI105 : in  std_logic;
    EI106 : in  std_logic;
    EI107 : in  std_logic;
    EI108 : in  std_logic;
    EI109 : in  std_logic;
    EI110 : in  std_logic;
    EI111 : in  std_logic;
    EI112 : in  std_logic;
    EI113 : in  std_logic;
    EI114 : in  std_logic;
    EI115 : in  std_logic;
    EI116 : in  std_logic;
    EI117 : in  std_logic;
    EI118 : in  std_logic;
    EI119 : in  std_logic;
    EI120 : in  std_logic;
    EI121 : in  std_logic;
    EI122 : in  std_logic;
    EI123 : in  std_logic;
    EI124 : in  std_logic;
    EI125 : in  std_logic;
    EI126 : in  std_logic;
    EI127 : in  std_logic;
    EI128 : in  std_logic;
    EI129 : in  std_logic;
    EI130 : in  std_logic;
    EI131 : in  std_logic;
    EI132 : in  std_logic;
    EI133 : in  std_logic;
    EI134 : in  std_logic;
    EI135 : in  std_logic;
    EI136 : in  std_logic;
    EI137 : in  std_logic;
    EI138 : in  std_logic;
    EI139 : in  std_logic;
    EI140 : in  std_logic;
    EI141 : in  std_logic;
    EI142 : in  std_logic;
    EI143 : in  std_logic;
    EI144 : in  std_logic;
    EI145 : in  std_logic;
    EI146 : in  std_logic;
    EI147 : in  std_logic;
    EI148 : in  std_logic;
    EI149 : in  std_logic;
    EI150 : in  std_logic;
    EI151 : in  std_logic;
    EI152 : in  std_logic;
    EI153 : in  std_logic;
    EI154 : in  std_logic;
    EI155 : in  std_logic;
    EI156 : in  std_logic;
    EI157 : in  std_logic;
    EI158 : in  std_logic;
    EI159 : in  std_logic;
    EI160 : in  std_logic;
    EI161 : in  std_logic;
    EI162 : in  std_logic;
    EI163 : in  std_logic;
    EI164 : in  std_logic;
    EI165 : in  std_logic;
    EI166 : in  std_logic;
    EI167 : in  std_logic;
    EI168 : in  std_logic;
    EI169 : in  std_logic;
    EI170 : in  std_logic;
    EI171 : in  std_logic;
    EI172 : in  std_logic;
    EI173 : in  std_logic;
    EI174 : in  std_logic;
    EI175 : in  std_logic;
    EI176 : in  std_logic;
    EI177 : in  std_logic;
    EI178 : in  std_logic;
    EI179 : in  std_logic;
    EI180 : in  std_logic;
    EI181 : in  std_logic;
    EI182 : in  std_logic;
    EI183 : in  std_logic;
    EI184 : in  std_logic;
    EI185 : in  std_logic;
    EI186 : in  std_logic;
    EI187 : in  std_logic;
    EI188 : in  std_logic;
    EI189 : in  std_logic;
    EI190 : in  std_logic;
    EI191 : in  std_logic;
    EI192 : in  std_logic;
    EI_CK : out std_logic;
    EO_CK : out std_logic;
    EO1   : out std_logic;
    EO2   : out std_logic;
    EO3   : out std_logic;
    EO4   : out std_logic;
    EO5   : out std_logic;
    EO6   : out std_logic;
    EO7   : out std_logic;
    EO8   : out std_logic;
    EO9   : out std_logic;
    EO10  : out std_logic;
    EO11  : out std_logic;
    EO12  : out std_logic;
    EO13  : out std_logic;
    EO14  : out std_logic;
    EO15  : out std_logic;
    EO16  : out std_logic;
    EO17  : out std_logic;
    EO18  : out std_logic;
    EO19  : out std_logic;
    EO20  : out std_logic;
    EO21  : out std_logic;
    EO22  : out std_logic;
    EO23  : out std_logic;
    EO24  : out std_logic;
    EO25  : out std_logic;
    EO26  : out std_logic;
    EO27  : out std_logic;
    EO28  : out std_logic;
    EO29  : out std_logic;
    EO30  : out std_logic;
    EO31  : out std_logic;
    EO32  : out std_logic;
    EO33  : out std_logic;
    EO34  : out std_logic;
    EO35  : out std_logic;
    EO36  : out std_logic;
    EO37  : out std_logic;
    EO38  : out std_logic;
    EO39  : out std_logic;
    EO40  : out std_logic;
    EO41  : out std_logic;
    EO42  : out std_logic;
    EO43  : out std_logic;
    EO44  : out std_logic;
    EO45  : out std_logic;
    EO46  : out std_logic;
    EO47  : out std_logic;
    EO48  : out std_logic;
    EO49  : out std_logic;
    EO50  : out std_logic;
    EO51  : out std_logic;
    EO52  : out std_logic;
    EO53  : out std_logic;
    EO54  : out std_logic;
    EO55  : out std_logic;
    EO56  : out std_logic;
    EO57  : out std_logic;
    EO58  : out std_logic;
    EO59  : out std_logic;
    EO60  : out std_logic;
    EO61  : out std_logic;
    EO62  : out std_logic;
    EO63  : out std_logic;
    EO64  : out std_logic;
    EO65  : out std_logic;
    EO66  : out std_logic;
    EO67  : out std_logic;
    EO68  : out std_logic;
    EO69  : out std_logic;
    EO70  : out std_logic;
    EO71  : out std_logic;
    EO72  : out std_logic;
    EO73  : out std_logic;
    EO74  : out std_logic;
    EO75  : out std_logic;
    EO76  : out std_logic;
    EO77  : out std_logic;
    EO78  : out std_logic;
    EO79  : out std_logic;
    EO80  : out std_logic;
    EO81  : out std_logic;
    EO82  : out std_logic;
    EO83  : out std_logic;
    EO84  : out std_logic;
    EO85  : out std_logic;
    EO86  : out std_logic;
    EO87  : out std_logic;
    EO88  : out std_logic;
    EO89  : out std_logic;
    EO90  : out std_logic;
    EO91  : out std_logic;
    EO92  : out std_logic;
    EO93  : out std_logic;
    EO94  : out std_logic;
    EO95  : out std_logic;
    EO96  : out std_logic;
    EO97  : out std_logic;
    EO98  : out std_logic;
    EO99  : out std_logic;
    EO100 : out std_logic;
    EO101 : out std_logic;
    EO102 : out std_logic;
    EO103 : out std_logic;
    EO104 : out std_logic;
    EO105 : out std_logic;
    EO106 : out std_logic;
    EO107 : out std_logic;
    EO108 : out std_logic;
    EO109 : out std_logic;
    EO110 : out std_logic;
    EO111 : out std_logic;
    EO112 : out std_logic;
    EO113 : out std_logic;
    EO114 : out std_logic;
    EO115 : out std_logic;
    EO116 : out std_logic;
    EO117 : out std_logic;
    EO118 : out std_logic;
    EO119 : out std_logic;
    EO120 : out std_logic;
    EO121 : out std_logic;
    EO122 : out std_logic;
    EO123 : out std_logic;
    EO124 : out std_logic;
    EO125 : out std_logic;
    EO126 : out std_logic;
    EO127 : out std_logic;
    EO128 : out std_logic;
    EO129 : out std_logic;
    EO130 : out std_logic;
    EO131 : out std_logic;
    EO132 : out std_logic;
    EO133 : out std_logic;
    EO134 : out std_logic;
    EO135 : out std_logic;
    EO136 : out std_logic;
    EO137 : out std_logic;
    EO138 : out std_logic;
    EO139 : out std_logic;
    EO140 : out std_logic;
    EO141 : out std_logic;
    EO142 : out std_logic;
    EO143 : out std_logic;
    EO144 : out std_logic;
    EO145 : out std_logic;
    EO146 : out std_logic;
    EO147 : out std_logic;
    EO148 : out std_logic;
    EO149 : out std_logic;
    EO150 : out std_logic;
    EO151 : out std_logic;
    EO152 : out std_logic;
    EO153 : out std_logic;
    EO154 : out std_logic;
    EO155 : out std_logic;
    EO156 : out std_logic;
    EO157 : out std_logic;
    EO158 : out std_logic;
    EO159 : out std_logic;
    EO160 : out std_logic;
    EO161 : out std_logic;
    EO162 : out std_logic;
    EO163 : out std_logic;
    EO164 : out std_logic;
    EO165 : out std_logic;
    EO166 : out std_logic;
    EO167 : out std_logic;
    EO168 : out std_logic;
    EO169 : out std_logic;
    EO170 : out std_logic;
    EO171 : out std_logic;
    EO172 : out std_logic;
    EO173 : out std_logic;
    EO174 : out std_logic;
    EO175 : out std_logic;
    EO176 : out std_logic;
    EO177 : out std_logic;
    EO178 : out std_logic;
    EO179 : out std_logic;
    EO180 : out std_logic;
    EO181 : out std_logic;
    EO182 : out std_logic;
    EO183 : out std_logic;
    EO184 : out std_logic;
    EO185 : out std_logic;
    EO186 : out std_logic;
    EO187 : out std_logic;
    EO188 : out std_logic;
    EO189 : out std_logic;
    EO190 : out std_logic;
    EO191 : out std_logic;
    EO192 : out std_logic;
    FI1   : in  std_logic;
    FI2   : in  std_logic;
    FI3   : in  std_logic;
    FI4   : in  std_logic;
    FI5   : in  std_logic;
    FI6   : in  std_logic;
    FI7   : in  std_logic;
    FI8   : in  std_logic;
    FI9   : in  std_logic;
    FI10  : in  std_logic;
    FI11  : in  std_logic;
    FI12  : in  std_logic;
    FI13  : in  std_logic;
    FI14  : in  std_logic;
    FI15  : in  std_logic;
    FI16  : in  std_logic;
    FI17  : in  std_logic;
    FI18  : in  std_logic;
    FI19  : in  std_logic;
    FI20  : in  std_logic;
    FI21  : in  std_logic;
    FI22  : in  std_logic;
    FI23  : in  std_logic;
    FI24  : in  std_logic;
    FI25  : in  std_logic;
    FI26  : in  std_logic;
    FI27  : in  std_logic;
    FI28  : in  std_logic;
    FI29  : in  std_logic;
    FI30  : in  std_logic;
    FI31  : in  std_logic;
    FI32  : in  std_logic;
    FI33  : in  std_logic;
    FI34  : in  std_logic;
    FI35  : in  std_logic;
    FI36  : in  std_logic;
    FI37  : in  std_logic;
    FI38  : in  std_logic;
    FI39  : in  std_logic;
    FI40  : in  std_logic;
    FI41  : in  std_logic;
    FI42  : in  std_logic;
    FI43  : in  std_logic;
    FI44  : in  std_logic;
    FI45  : in  std_logic;
    FI46  : in  std_logic;
    FI47  : in  std_logic;
    FI48  : in  std_logic;
    FI49  : in  std_logic;
    FI50  : in  std_logic;
    FI51  : in  std_logic;
    FI52  : in  std_logic;
    FI53  : in  std_logic;
    FI54  : in  std_logic;
    FI55  : in  std_logic;
    FI56  : in  std_logic;
    FI57  : in  std_logic;
    FI58  : in  std_logic;
    FI59  : in  std_logic;
    FI60  : in  std_logic;
    FI61  : in  std_logic;
    FI62  : in  std_logic;
    FI63  : in  std_logic;
    FI64  : in  std_logic;
    FI65  : in  std_logic;
    FI66  : in  std_logic;
    FI67  : in  std_logic;
    FI68  : in  std_logic;
    FI69  : in  std_logic;
    FI70  : in  std_logic;
    FI71  : in  std_logic;
    FI72  : in  std_logic;
    FI73  : in  std_logic;
    FI74  : in  std_logic;
    FI75  : in  std_logic;
    FI76  : in  std_logic;
    FI77  : in  std_logic;
    FI78  : in  std_logic;
    FI79  : in  std_logic;
    FI80  : in  std_logic;
    FI81  : in  std_logic;
    FI82  : in  std_logic;
    FI83  : in  std_logic;
    FI84  : in  std_logic;
    FI85  : in  std_logic;
    FI86  : in  std_logic;
    FI87  : in  std_logic;
    FI88  : in  std_logic;
    FI89  : in  std_logic;
    FI90  : in  std_logic;
    FI91  : in  std_logic;
    FI92  : in  std_logic;
    FI93  : in  std_logic;
    FI94  : in  std_logic;
    FI95  : in  std_logic;
    FI96  : in  std_logic;
    FI97  : in  std_logic;
    FI98  : in  std_logic;
    FI99  : in  std_logic;
    FI100 : in  std_logic;
    FI101 : in  std_logic;
    FI102 : in  std_logic;
    FI103 : in  std_logic;
    FI104 : in  std_logic;
    FI105 : in  std_logic;
    FI106 : in  std_logic;
    FI107 : in  std_logic;
    FI108 : in  std_logic;
    FI109 : in  std_logic;
    FI110 : in  std_logic;
    FI111 : in  std_logic;
    FI112 : in  std_logic;
    FI113 : in  std_logic;
    FI114 : in  std_logic;
    FI115 : in  std_logic;
    FI116 : in  std_logic;
    FI117 : in  std_logic;
    FI118 : in  std_logic;
    FI119 : in  std_logic;
    FI120 : in  std_logic;
    FI121 : in  std_logic;
    FI122 : in  std_logic;
    FI123 : in  std_logic;
    FI124 : in  std_logic;
    FI125 : in  std_logic;
    FI126 : in  std_logic;
    FI127 : in  std_logic;
    FI128 : in  std_logic;
    FI129 : in  std_logic;
    FI130 : in  std_logic;
    FI131 : in  std_logic;
    FI132 : in  std_logic;
    FI133 : in  std_logic;
    FI134 : in  std_logic;
    FI135 : in  std_logic;
    FI136 : in  std_logic;
    FI137 : in  std_logic;
    FI138 : in  std_logic;
    FI139 : in  std_logic;
    FI140 : in  std_logic;
    FI141 : in  std_logic;
    FI142 : in  std_logic;
    FI143 : in  std_logic;
    FI144 : in  std_logic;
    FI145 : in  std_logic;
    FI146 : in  std_logic;
    FI147 : in  std_logic;
    FI148 : in  std_logic;
    FI149 : in  std_logic;
    FI150 : in  std_logic;
    FI151 : in  std_logic;
    FI152 : in  std_logic;
    FI153 : in  std_logic;
    FI154 : in  std_logic;
    FI155 : in  std_logic;
    FI156 : in  std_logic;
    FI157 : in  std_logic;
    FI158 : in  std_logic;
    FI159 : in  std_logic;
    FI160 : in  std_logic;
    FI161 : in  std_logic;
    FI162 : in  std_logic;
    FI163 : in  std_logic;
    FI164 : in  std_logic;
    FI165 : in  std_logic;
    FI166 : in  std_logic;
    FI167 : in  std_logic;
    FI168 : in  std_logic;
    FI169 : in  std_logic;
    FI170 : in  std_logic;
    FI171 : in  std_logic;
    FI172 : in  std_logic;
    FI173 : in  std_logic;
    FI174 : in  std_logic;
    FI175 : in  std_logic;
    FI176 : in  std_logic;
    FI177 : in  std_logic;
    FI178 : in  std_logic;
    FI179 : in  std_logic;
    FI180 : in  std_logic;
    FI181 : in  std_logic;
    FI182 : in  std_logic;
    FI183 : in  std_logic;
    FI184 : in  std_logic;
    FI185 : in  std_logic;
    FI186 : in  std_logic;
    FI187 : in  std_logic;
    FI188 : in  std_logic;
    FI189 : in  std_logic;
    FI190 : in  std_logic;
    FI191 : in  std_logic;
    FI192 : in  std_logic;
    FO1   : out std_logic;
    FO2   : out std_logic;
    FO3   : out std_logic;
    FO4   : out std_logic;
    FO5   : out std_logic;
    FO6   : out std_logic;
    FO7   : out std_logic;
    FO8   : out std_logic;
    FO9   : out std_logic;
    FO10  : out std_logic;
    FO11  : out std_logic;
    FO12  : out std_logic;
    FO13  : out std_logic;
    FO14  : out std_logic;
    FO15  : out std_logic;
    FO16  : out std_logic;
    FO17  : out std_logic;
    FO18  : out std_logic;
    FO19  : out std_logic;
    FO20  : out std_logic;
    FO21  : out std_logic;
    FO22  : out std_logic;
    FO23  : out std_logic;
    FO24  : out std_logic;
    FO25  : out std_logic;
    FO26  : out std_logic;
    FO27  : out std_logic;
    FO28  : out std_logic;
    FO29  : out std_logic;
    FO30  : out std_logic;
    FO31  : out std_logic;
    FO32  : out std_logic;
    FO33  : out std_logic;
    FO34  : out std_logic;
    FO35  : out std_logic;
    FO36  : out std_logic;
    FO37  : out std_logic;
    FO38  : out std_logic;
    FO39  : out std_logic;
    FO40  : out std_logic;
    FO41  : out std_logic;
    FO42  : out std_logic;
    FO43  : out std_logic;
    FO44  : out std_logic;
    FO45  : out std_logic;
    FO46  : out std_logic;
    FO47  : out std_logic;
    FO48  : out std_logic;
    FO49  : out std_logic;
    FO50  : out std_logic;
    FO51  : out std_logic;
    FO52  : out std_logic;
    FO53  : out std_logic;
    FO54  : out std_logic;
    FO55  : out std_logic;
    FO56  : out std_logic;
    FO57  : out std_logic;
    FO58  : out std_logic;
    FO59  : out std_logic;
    FO60  : out std_logic;
    FO61  : out std_logic;
    FO62  : out std_logic;
    FO63  : out std_logic;
    FO64  : out std_logic;
    FO65  : out std_logic;
    FO66  : out std_logic;
    FO67  : out std_logic;
    FO68  : out std_logic;
    FO69  : out std_logic;
    FO70  : out std_logic;
    FO71  : out std_logic;
    FO72  : out std_logic;
    FO73  : out std_logic;
    FO74  : out std_logic;
    FO75  : out std_logic;
    FO76  : out std_logic;
    FO77  : out std_logic;
    FO78  : out std_logic;
    FO79  : out std_logic;
    FO80  : out std_logic;
    FO81  : out std_logic;
    FO82  : out std_logic;
    FO83  : out std_logic;
    FO84  : out std_logic;
    FO85  : out std_logic;
    FO86  : out std_logic;
    FO87  : out std_logic;
    FO88  : out std_logic;
    FO89  : out std_logic;
    FO90  : out std_logic;
    FO91  : out std_logic;
    FO92  : out std_logic;
    FO93  : out std_logic;
    FO94  : out std_logic;
    FO95  : out std_logic;
    FO96  : out std_logic;
    FO97  : out std_logic;
    FO98  : out std_logic;
    FO99  : out std_logic;
    FO100 : out std_logic;
    FO101 : out std_logic;
    FO102 : out std_logic;
    FO103 : out std_logic;
    FO104 : out std_logic;
    FO105 : out std_logic;
    FO106 : out std_logic;
    FO107 : out std_logic;
    FO108 : out std_logic;
    FO109 : out std_logic;
    FO110 : out std_logic;
    FO111 : out std_logic;
    FO112 : out std_logic;
    FO113 : out std_logic;
    FO114 : out std_logic;
    FO115 : out std_logic;
    FO116 : out std_logic;
    FO117 : out std_logic;
    FO118 : out std_logic;
    FO119 : out std_logic;
    FO120 : out std_logic;
    FO121 : out std_logic;
    FO122 : out std_logic;
    FO123 : out std_logic;
    FO124 : out std_logic;
    FO125 : out std_logic;
    FO126 : out std_logic;
    FO127 : out std_logic;
    FO128 : out std_logic;
    FO129 : out std_logic;
    FO130 : out std_logic;
    FO131 : out std_logic;
    FO132 : out std_logic;
    FO133 : out std_logic;
    FO134 : out std_logic;
    FO135 : out std_logic;
    FO136 : out std_logic;
    FO137 : out std_logic;
    FO138 : out std_logic;
    FO139 : out std_logic;
    FO140 : out std_logic;
    FO141 : out std_logic;
    FO142 : out std_logic;
    FO143 : out std_logic;
    FO144 : out std_logic;
    FO145 : out std_logic;
    FO146 : out std_logic;
    FO147 : out std_logic;
    FO148 : out std_logic;
    FO149 : out std_logic;
    FO150 : out std_logic;
    FO151 : out std_logic;
    FO152 : out std_logic;
    FO153 : out std_logic;
    FO154 : out std_logic;
    FO155 : out std_logic;
    FO156 : out std_logic;
    FO157 : out std_logic;
    FO158 : out std_logic;
    FO159 : out std_logic;
    FO160 : out std_logic;
    FO161 : out std_logic;
    FO162 : out std_logic;
    FO163 : out std_logic;
    FO164 : out std_logic;
    FO165 : out std_logic;
    FO166 : out std_logic;
    FO167 : out std_logic;
    FO168 : out std_logic;
    FO169 : out std_logic;
    FO170 : out std_logic;
    FO171 : out std_logic;
    FO172 : out std_logic;
    FO173 : out std_logic;
    FO174 : out std_logic;
    FO175 : out std_logic;
    FO176 : out std_logic;
    FO177 : out std_logic;
    FO178 : out std_logic;
    FO179 : out std_logic;
    FO180 : out std_logic;
    FO181 : out std_logic;
    FO182 : out std_logic;
    FO183 : out std_logic;
    FO184 : out std_logic;
    FO185 : out std_logic;
    FO186 : out std_logic;
    FO187 : out std_logic;
    FO188 : out std_logic;
    FO189 : out std_logic;
    FO190 : out std_logic;
    FO191 : out std_logic;
    FO192 : out std_logic
);
end NX_RB;

architecture NX_RTL of NX_RB is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RB";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RB_WRAP definition                                                              2017/06/18
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_RB_WRAP is
generic (
    -- input : EI to FO
    inputClk      : bit_vector( 1 downto 0) := B"00"; -- 00 = CK[0], 01 = CK[1], 10 = CK[2] and 11 = CK[3]
    inputBypass   : bit_vector(23 downto 0) := B"000000000000000000000000"; -- 1 bypass active, LSB is bypass registers 0 to 7 ... MSB is bypass registers 183 to 191
    -- output : FI to EO
    inputContext  : string := ""; -- input context intialization
    outputClk     : bit_vector( 1 downto 0) := B"00"; -- 00 = CK[0], 01 = CK[1], 10 = CK[2] and 11 = CK[3]
    outputBypass  : bit_vector(23 downto 0) := B"000000000000000000000000";  -- 1 bypass active, LSB is bypass registers 1 to 8 ... MSB is bypass registers 184 to 192
    outputContext : string := "" -- output context intialization
);
port (
    CK      : in  std_logic_vector(  3 downto 0);
    EI_CK   : out std_logic;
    EO_CK   : out std_logic;
    EI      : in  std_logic_vector(191 downto 0);
    EO      : out std_logic_vector(191 downto 0);
    FI      : in  std_logic_vector(191 downto 0);
    FO      : out std_logic_vector(191 downto 0)
);
end NX_RB_WRAP;

architecture NX_RTL of NX_RB_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RB
generic (
    inputClk      : bit_vector( 1 downto 0) := B"00";
    inputBypass   : bit_vector(23 downto 0) := B"000000000000000000000000";
    inputContext  : string := "";
    outputClk     : bit_vector( 1 downto 0) := B"00";
    outputBypass  : bit_vector(23 downto 0) := B"000000000000000000000000";
    outputContext : string := ""
);
port (
    CK1   : in  std_logic;
    CK2   : in  std_logic;
    CK3   : in  std_logic;
    CK4   : in  std_logic;
    EI1   : in  std_logic;
    EI2   : in  std_logic;
    EI3   : in  std_logic;
    EI4   : in  std_logic;
    EI5   : in  std_logic;
    EI6   : in  std_logic;
    EI7   : in  std_logic;
    EI8   : in  std_logic;
    EI9   : in  std_logic;
    EI10  : in  std_logic;
    EI11  : in  std_logic;
    EI12  : in  std_logic;
    EI13  : in  std_logic;
    EI14  : in  std_logic;
    EI15  : in  std_logic;
    EI16  : in  std_logic;
    EI17  : in  std_logic;
    EI18  : in  std_logic;
    EI19  : in  std_logic;
    EI20  : in  std_logic;
    EI21  : in  std_logic;
    EI22  : in  std_logic;
    EI23  : in  std_logic;
    EI24  : in  std_logic;
    EI25  : in  std_logic;
    EI26  : in  std_logic;
    EI27  : in  std_logic;
    EI28  : in  std_logic;
    EI29  : in  std_logic;
    EI30  : in  std_logic;
    EI31  : in  std_logic;
    EI32  : in  std_logic;
    EI33  : in  std_logic;
    EI34  : in  std_logic;
    EI35  : in  std_logic;
    EI36  : in  std_logic;
    EI37  : in  std_logic;
    EI38  : in  std_logic;
    EI39  : in  std_logic;
    EI40  : in  std_logic;
    EI41  : in  std_logic;
    EI42  : in  std_logic;
    EI43  : in  std_logic;
    EI44  : in  std_logic;
    EI45  : in  std_logic;
    EI46  : in  std_logic;
    EI47  : in  std_logic;
    EI48  : in  std_logic;
    EI49  : in  std_logic;
    EI50  : in  std_logic;
    EI51  : in  std_logic;
    EI52  : in  std_logic;
    EI53  : in  std_logic;
    EI54  : in  std_logic;
    EI55  : in  std_logic;
    EI56  : in  std_logic;
    EI57  : in  std_logic;
    EI58  : in  std_logic;
    EI59  : in  std_logic;
    EI60  : in  std_logic;
    EI61  : in  std_logic;
    EI62  : in  std_logic;
    EI63  : in  std_logic;
    EI64  : in  std_logic;
    EI65  : in  std_logic;
    EI66  : in  std_logic;
    EI67  : in  std_logic;
    EI68  : in  std_logic;
    EI69  : in  std_logic;
    EI70  : in  std_logic;
    EI71  : in  std_logic;
    EI72  : in  std_logic;
    EI73  : in  std_logic;
    EI74  : in  std_logic;
    EI75  : in  std_logic;
    EI76  : in  std_logic;
    EI77  : in  std_logic;
    EI78  : in  std_logic;
    EI79  : in  std_logic;
    EI80  : in  std_logic;
    EI81  : in  std_logic;
    EI82  : in  std_logic;
    EI83  : in  std_logic;
    EI84  : in  std_logic;
    EI85  : in  std_logic;
    EI86  : in  std_logic;
    EI87  : in  std_logic;
    EI88  : in  std_logic;
    EI89  : in  std_logic;
    EI90  : in  std_logic;
    EI91  : in  std_logic;
    EI92  : in  std_logic;
    EI93  : in  std_logic;
    EI94  : in  std_logic;
    EI95  : in  std_logic;
    EI96  : in  std_logic;
    EI97  : in  std_logic;
    EI98  : in  std_logic;
    EI99  : in  std_logic;
    EI100 : in  std_logic;
    EI101 : in  std_logic;
    EI102 : in  std_logic;
    EI103 : in  std_logic;
    EI104 : in  std_logic;
    EI105 : in  std_logic;
    EI106 : in  std_logic;
    EI107 : in  std_logic;
    EI108 : in  std_logic;
    EI109 : in  std_logic;
    EI110 : in  std_logic;
    EI111 : in  std_logic;
    EI112 : in  std_logic;
    EI113 : in  std_logic;
    EI114 : in  std_logic;
    EI115 : in  std_logic;
    EI116 : in  std_logic;
    EI117 : in  std_logic;
    EI118 : in  std_logic;
    EI119 : in  std_logic;
    EI120 : in  std_logic;
    EI121 : in  std_logic;
    EI122 : in  std_logic;
    EI123 : in  std_logic;
    EI124 : in  std_logic;
    EI125 : in  std_logic;
    EI126 : in  std_logic;
    EI127 : in  std_logic;
    EI128 : in  std_logic;
    EI129 : in  std_logic;
    EI130 : in  std_logic;
    EI131 : in  std_logic;
    EI132 : in  std_logic;
    EI133 : in  std_logic;
    EI134 : in  std_logic;
    EI135 : in  std_logic;
    EI136 : in  std_logic;
    EI137 : in  std_logic;
    EI138 : in  std_logic;
    EI139 : in  std_logic;
    EI140 : in  std_logic;
    EI141 : in  std_logic;
    EI142 : in  std_logic;
    EI143 : in  std_logic;
    EI144 : in  std_logic;
    EI145 : in  std_logic;
    EI146 : in  std_logic;
    EI147 : in  std_logic;
    EI148 : in  std_logic;
    EI149 : in  std_logic;
    EI150 : in  std_logic;
    EI151 : in  std_logic;
    EI152 : in  std_logic;
    EI153 : in  std_logic;
    EI154 : in  std_logic;
    EI155 : in  std_logic;
    EI156 : in  std_logic;
    EI157 : in  std_logic;
    EI158 : in  std_logic;
    EI159 : in  std_logic;
    EI160 : in  std_logic;
    EI161 : in  std_logic;
    EI162 : in  std_logic;
    EI163 : in  std_logic;
    EI164 : in  std_logic;
    EI165 : in  std_logic;
    EI166 : in  std_logic;
    EI167 : in  std_logic;
    EI168 : in  std_logic;
    EI169 : in  std_logic;
    EI170 : in  std_logic;
    EI171 : in  std_logic;
    EI172 : in  std_logic;
    EI173 : in  std_logic;
    EI174 : in  std_logic;
    EI175 : in  std_logic;
    EI176 : in  std_logic;
    EI177 : in  std_logic;
    EI178 : in  std_logic;
    EI179 : in  std_logic;
    EI180 : in  std_logic;
    EI181 : in  std_logic;
    EI182 : in  std_logic;
    EI183 : in  std_logic;
    EI184 : in  std_logic;
    EI185 : in  std_logic;
    EI186 : in  std_logic;
    EI187 : in  std_logic;
    EI188 : in  std_logic;
    EI189 : in  std_logic;
    EI190 : in  std_logic;
    EI191 : in  std_logic;
    EI192 : in  std_logic;
    EI_CK : out std_logic;
    EO_CK : out std_logic;
    EO1   : out std_logic;
    EO2   : out std_logic;
    EO3   : out std_logic;
    EO4   : out std_logic;
    EO5   : out std_logic;
    EO6   : out std_logic;
    EO7   : out std_logic;
    EO8   : out std_logic;
    EO9   : out std_logic;
    EO10  : out std_logic;
    EO11  : out std_logic;
    EO12  : out std_logic;
    EO13  : out std_logic;
    EO14  : out std_logic;
    EO15  : out std_logic;
    EO16  : out std_logic;
    EO17  : out std_logic;
    EO18  : out std_logic;
    EO19  : out std_logic;
    EO20  : out std_logic;
    EO21  : out std_logic;
    EO22  : out std_logic;
    EO23  : out std_logic;
    EO24  : out std_logic;
    EO25  : out std_logic;
    EO26  : out std_logic;
    EO27  : out std_logic;
    EO28  : out std_logic;
    EO29  : out std_logic;
    EO30  : out std_logic;
    EO31  : out std_logic;
    EO32  : out std_logic;
    EO33  : out std_logic;
    EO34  : out std_logic;
    EO35  : out std_logic;
    EO36  : out std_logic;
    EO37  : out std_logic;
    EO38  : out std_logic;
    EO39  : out std_logic;
    EO40  : out std_logic;
    EO41  : out std_logic;
    EO42  : out std_logic;
    EO43  : out std_logic;
    EO44  : out std_logic;
    EO45  : out std_logic;
    EO46  : out std_logic;
    EO47  : out std_logic;
    EO48  : out std_logic;
    EO49  : out std_logic;
    EO50  : out std_logic;
    EO51  : out std_logic;
    EO52  : out std_logic;
    EO53  : out std_logic;
    EO54  : out std_logic;
    EO55  : out std_logic;
    EO56  : out std_logic;
    EO57  : out std_logic;
    EO58  : out std_logic;
    EO59  : out std_logic;
    EO60  : out std_logic;
    EO61  : out std_logic;
    EO62  : out std_logic;
    EO63  : out std_logic;
    EO64  : out std_logic;
    EO65  : out std_logic;
    EO66  : out std_logic;
    EO67  : out std_logic;
    EO68  : out std_logic;
    EO69  : out std_logic;
    EO70  : out std_logic;
    EO71  : out std_logic;
    EO72  : out std_logic;
    EO73  : out std_logic;
    EO74  : out std_logic;
    EO75  : out std_logic;
    EO76  : out std_logic;
    EO77  : out std_logic;
    EO78  : out std_logic;
    EO79  : out std_logic;
    EO80  : out std_logic;
    EO81  : out std_logic;
    EO82  : out std_logic;
    EO83  : out std_logic;
    EO84  : out std_logic;
    EO85  : out std_logic;
    EO86  : out std_logic;
    EO87  : out std_logic;
    EO88  : out std_logic;
    EO89  : out std_logic;
    EO90  : out std_logic;
    EO91  : out std_logic;
    EO92  : out std_logic;
    EO93  : out std_logic;
    EO94  : out std_logic;
    EO95  : out std_logic;
    EO96  : out std_logic;
    EO97  : out std_logic;
    EO98  : out std_logic;
    EO99  : out std_logic;
    EO100 : out std_logic;
    EO101 : out std_logic;
    EO102 : out std_logic;
    EO103 : out std_logic;
    EO104 : out std_logic;
    EO105 : out std_logic;
    EO106 : out std_logic;
    EO107 : out std_logic;
    EO108 : out std_logic;
    EO109 : out std_logic;
    EO110 : out std_logic;
    EO111 : out std_logic;
    EO112 : out std_logic;
    EO113 : out std_logic;
    EO114 : out std_logic;
    EO115 : out std_logic;
    EO116 : out std_logic;
    EO117 : out std_logic;
    EO118 : out std_logic;
    EO119 : out std_logic;
    EO120 : out std_logic;
    EO121 : out std_logic;
    EO122 : out std_logic;
    EO123 : out std_logic;
    EO124 : out std_logic;
    EO125 : out std_logic;
    EO126 : out std_logic;
    EO127 : out std_logic;
    EO128 : out std_logic;
    EO129 : out std_logic;
    EO130 : out std_logic;
    EO131 : out std_logic;
    EO132 : out std_logic;
    EO133 : out std_logic;
    EO134 : out std_logic;
    EO135 : out std_logic;
    EO136 : out std_logic;
    EO137 : out std_logic;
    EO138 : out std_logic;
    EO139 : out std_logic;
    EO140 : out std_logic;
    EO141 : out std_logic;
    EO142 : out std_logic;
    EO143 : out std_logic;
    EO144 : out std_logic;
    EO145 : out std_logic;
    EO146 : out std_logic;
    EO147 : out std_logic;
    EO148 : out std_logic;
    EO149 : out std_logic;
    EO150 : out std_logic;
    EO151 : out std_logic;
    EO152 : out std_logic;
    EO153 : out std_logic;
    EO154 : out std_logic;
    EO155 : out std_logic;
    EO156 : out std_logic;
    EO157 : out std_logic;
    EO158 : out std_logic;
    EO159 : out std_logic;
    EO160 : out std_logic;
    EO161 : out std_logic;
    EO162 : out std_logic;
    EO163 : out std_logic;
    EO164 : out std_logic;
    EO165 : out std_logic;
    EO166 : out std_logic;
    EO167 : out std_logic;
    EO168 : out std_logic;
    EO169 : out std_logic;
    EO170 : out std_logic;
    EO171 : out std_logic;
    EO172 : out std_logic;
    EO173 : out std_logic;
    EO174 : out std_logic;
    EO175 : out std_logic;
    EO176 : out std_logic;
    EO177 : out std_logic;
    EO178 : out std_logic;
    EO179 : out std_logic;
    EO180 : out std_logic;
    EO181 : out std_logic;
    EO182 : out std_logic;
    EO183 : out std_logic;
    EO184 : out std_logic;
    EO185 : out std_logic;
    EO186 : out std_logic;
    EO187 : out std_logic;
    EO188 : out std_logic;
    EO189 : out std_logic;
    EO190 : out std_logic;
    EO191 : out std_logic;
    EO192 : out std_logic;
    FI1   : in  std_logic;
    FI2   : in  std_logic;
    FI3   : in  std_logic;
    FI4   : in  std_logic;
    FI5   : in  std_logic;
    FI6   : in  std_logic;
    FI7   : in  std_logic;
    FI8   : in  std_logic;
    FI9   : in  std_logic;
    FI10  : in  std_logic;
    FI11  : in  std_logic;
    FI12  : in  std_logic;
    FI13  : in  std_logic;
    FI14  : in  std_logic;
    FI15  : in  std_logic;
    FI16  : in  std_logic;
    FI17  : in  std_logic;
    FI18  : in  std_logic;
    FI19  : in  std_logic;
    FI20  : in  std_logic;
    FI21  : in  std_logic;
    FI22  : in  std_logic;
    FI23  : in  std_logic;
    FI24  : in  std_logic;
    FI25  : in  std_logic;
    FI26  : in  std_logic;
    FI27  : in  std_logic;
    FI28  : in  std_logic;
    FI29  : in  std_logic;
    FI30  : in  std_logic;
    FI31  : in  std_logic;
    FI32  : in  std_logic;
    FI33  : in  std_logic;
    FI34  : in  std_logic;
    FI35  : in  std_logic;
    FI36  : in  std_logic;
    FI37  : in  std_logic;
    FI38  : in  std_logic;
    FI39  : in  std_logic;
    FI40  : in  std_logic;
    FI41  : in  std_logic;
    FI42  : in  std_logic;
    FI43  : in  std_logic;
    FI44  : in  std_logic;
    FI45  : in  std_logic;
    FI46  : in  std_logic;
    FI47  : in  std_logic;
    FI48  : in  std_logic;
    FI49  : in  std_logic;
    FI50  : in  std_logic;
    FI51  : in  std_logic;
    FI52  : in  std_logic;
    FI53  : in  std_logic;
    FI54  : in  std_logic;
    FI55  : in  std_logic;
    FI56  : in  std_logic;
    FI57  : in  std_logic;
    FI58  : in  std_logic;
    FI59  : in  std_logic;
    FI60  : in  std_logic;
    FI61  : in  std_logic;
    FI62  : in  std_logic;
    FI63  : in  std_logic;
    FI64  : in  std_logic;
    FI65  : in  std_logic;
    FI66  : in  std_logic;
    FI67  : in  std_logic;
    FI68  : in  std_logic;
    FI69  : in  std_logic;
    FI70  : in  std_logic;
    FI71  : in  std_logic;
    FI72  : in  std_logic;
    FI73  : in  std_logic;
    FI74  : in  std_logic;
    FI75  : in  std_logic;
    FI76  : in  std_logic;
    FI77  : in  std_logic;
    FI78  : in  std_logic;
    FI79  : in  std_logic;
    FI80  : in  std_logic;
    FI81  : in  std_logic;
    FI82  : in  std_logic;
    FI83  : in  std_logic;
    FI84  : in  std_logic;
    FI85  : in  std_logic;
    FI86  : in  std_logic;
    FI87  : in  std_logic;
    FI88  : in  std_logic;
    FI89  : in  std_logic;
    FI90  : in  std_logic;
    FI91  : in  std_logic;
    FI92  : in  std_logic;
    FI93  : in  std_logic;
    FI94  : in  std_logic;
    FI95  : in  std_logic;
    FI96  : in  std_logic;
    FI97  : in  std_logic;
    FI98  : in  std_logic;
    FI99  : in  std_logic;
    FI100 : in  std_logic;
    FI101 : in  std_logic;
    FI102 : in  std_logic;
    FI103 : in  std_logic;
    FI104 : in  std_logic;
    FI105 : in  std_logic;
    FI106 : in  std_logic;
    FI107 : in  std_logic;
    FI108 : in  std_logic;
    FI109 : in  std_logic;
    FI110 : in  std_logic;
    FI111 : in  std_logic;
    FI112 : in  std_logic;
    FI113 : in  std_logic;
    FI114 : in  std_logic;
    FI115 : in  std_logic;
    FI116 : in  std_logic;
    FI117 : in  std_logic;
    FI118 : in  std_logic;
    FI119 : in  std_logic;
    FI120 : in  std_logic;
    FI121 : in  std_logic;
    FI122 : in  std_logic;
    FI123 : in  std_logic;
    FI124 : in  std_logic;
    FI125 : in  std_logic;
    FI126 : in  std_logic;
    FI127 : in  std_logic;
    FI128 : in  std_logic;
    FI129 : in  std_logic;
    FI130 : in  std_logic;
    FI131 : in  std_logic;
    FI132 : in  std_logic;
    FI133 : in  std_logic;
    FI134 : in  std_logic;
    FI135 : in  std_logic;
    FI136 : in  std_logic;
    FI137 : in  std_logic;
    FI138 : in  std_logic;
    FI139 : in  std_logic;
    FI140 : in  std_logic;
    FI141 : in  std_logic;
    FI142 : in  std_logic;
    FI143 : in  std_logic;
    FI144 : in  std_logic;
    FI145 : in  std_logic;
    FI146 : in  std_logic;
    FI147 : in  std_logic;
    FI148 : in  std_logic;
    FI149 : in  std_logic;
    FI150 : in  std_logic;
    FI151 : in  std_logic;
    FI152 : in  std_logic;
    FI153 : in  std_logic;
    FI154 : in  std_logic;
    FI155 : in  std_logic;
    FI156 : in  std_logic;
    FI157 : in  std_logic;
    FI158 : in  std_logic;
    FI159 : in  std_logic;
    FI160 : in  std_logic;
    FI161 : in  std_logic;
    FI162 : in  std_logic;
    FI163 : in  std_logic;
    FI164 : in  std_logic;
    FI165 : in  std_logic;
    FI166 : in  std_logic;
    FI167 : in  std_logic;
    FI168 : in  std_logic;
    FI169 : in  std_logic;
    FI170 : in  std_logic;
    FI171 : in  std_logic;
    FI172 : in  std_logic;
    FI173 : in  std_logic;
    FI174 : in  std_logic;
    FI175 : in  std_logic;
    FI176 : in  std_logic;
    FI177 : in  std_logic;
    FI178 : in  std_logic;
    FI179 : in  std_logic;
    FI180 : in  std_logic;
    FI181 : in  std_logic;
    FI182 : in  std_logic;
    FI183 : in  std_logic;
    FI184 : in  std_logic;
    FI185 : in  std_logic;
    FI186 : in  std_logic;
    FI187 : in  std_logic;
    FI188 : in  std_logic;
    FI189 : in  std_logic;
    FI190 : in  std_logic;
    FI191 : in  std_logic;
    FI192 : in  std_logic;
    FO1   : out std_logic;
    FO2   : out std_logic;
    FO3   : out std_logic;
    FO4   : out std_logic;
    FO5   : out std_logic;
    FO6   : out std_logic;
    FO7   : out std_logic;
    FO8   : out std_logic;
    FO9   : out std_logic;
    FO10  : out std_logic;
    FO11  : out std_logic;
    FO12  : out std_logic;
    FO13  : out std_logic;
    FO14  : out std_logic;
    FO15  : out std_logic;
    FO16  : out std_logic;
    FO17  : out std_logic;
    FO18  : out std_logic;
    FO19  : out std_logic;
    FO20  : out std_logic;
    FO21  : out std_logic;
    FO22  : out std_logic;
    FO23  : out std_logic;
    FO24  : out std_logic;
    FO25  : out std_logic;
    FO26  : out std_logic;
    FO27  : out std_logic;
    FO28  : out std_logic;
    FO29  : out std_logic;
    FO30  : out std_logic;
    FO31  : out std_logic;
    FO32  : out std_logic;
    FO33  : out std_logic;
    FO34  : out std_logic;
    FO35  : out std_logic;
    FO36  : out std_logic;
    FO37  : out std_logic;
    FO38  : out std_logic;
    FO39  : out std_logic;
    FO40  : out std_logic;
    FO41  : out std_logic;
    FO42  : out std_logic;
    FO43  : out std_logic;
    FO44  : out std_logic;
    FO45  : out std_logic;
    FO46  : out std_logic;
    FO47  : out std_logic;
    FO48  : out std_logic;
    FO49  : out std_logic;
    FO50  : out std_logic;
    FO51  : out std_logic;
    FO52  : out std_logic;
    FO53  : out std_logic;
    FO54  : out std_logic;
    FO55  : out std_logic;
    FO56  : out std_logic;
    FO57  : out std_logic;
    FO58  : out std_logic;
    FO59  : out std_logic;
    FO60  : out std_logic;
    FO61  : out std_logic;
    FO62  : out std_logic;
    FO63  : out std_logic;
    FO64  : out std_logic;
    FO65  : out std_logic;
    FO66  : out std_logic;
    FO67  : out std_logic;
    FO68  : out std_logic;
    FO69  : out std_logic;
    FO70  : out std_logic;
    FO71  : out std_logic;
    FO72  : out std_logic;
    FO73  : out std_logic;
    FO74  : out std_logic;
    FO75  : out std_logic;
    FO76  : out std_logic;
    FO77  : out std_logic;
    FO78  : out std_logic;
    FO79  : out std_logic;
    FO80  : out std_logic;
    FO81  : out std_logic;
    FO82  : out std_logic;
    FO83  : out std_logic;
    FO84  : out std_logic;
    FO85  : out std_logic;
    FO86  : out std_logic;
    FO87  : out std_logic;
    FO88  : out std_logic;
    FO89  : out std_logic;
    FO90  : out std_logic;
    FO91  : out std_logic;
    FO92  : out std_logic;
    FO93  : out std_logic;
    FO94  : out std_logic;
    FO95  : out std_logic;
    FO96  : out std_logic;
    FO97  : out std_logic;
    FO98  : out std_logic;
    FO99  : out std_logic;
    FO100 : out std_logic;
    FO101 : out std_logic;
    FO102 : out std_logic;
    FO103 : out std_logic;
    FO104 : out std_logic;
    FO105 : out std_logic;
    FO106 : out std_logic;
    FO107 : out std_logic;
    FO108 : out std_logic;
    FO109 : out std_logic;
    FO110 : out std_logic;
    FO111 : out std_logic;
    FO112 : out std_logic;
    FO113 : out std_logic;
    FO114 : out std_logic;
    FO115 : out std_logic;
    FO116 : out std_logic;
    FO117 : out std_logic;
    FO118 : out std_logic;
    FO119 : out std_logic;
    FO120 : out std_logic;
    FO121 : out std_logic;
    FO122 : out std_logic;
    FO123 : out std_logic;
    FO124 : out std_logic;
    FO125 : out std_logic;
    FO126 : out std_logic;
    FO127 : out std_logic;
    FO128 : out std_logic;
    FO129 : out std_logic;
    FO130 : out std_logic;
    FO131 : out std_logic;
    FO132 : out std_logic;
    FO133 : out std_logic;
    FO134 : out std_logic;
    FO135 : out std_logic;
    FO136 : out std_logic;
    FO137 : out std_logic;
    FO138 : out std_logic;
    FO139 : out std_logic;
    FO140 : out std_logic;
    FO141 : out std_logic;
    FO142 : out std_logic;
    FO143 : out std_logic;
    FO144 : out std_logic;
    FO145 : out std_logic;
    FO146 : out std_logic;
    FO147 : out std_logic;
    FO148 : out std_logic;
    FO149 : out std_logic;
    FO150 : out std_logic;
    FO151 : out std_logic;
    FO152 : out std_logic;
    FO153 : out std_logic;
    FO154 : out std_logic;
    FO155 : out std_logic;
    FO156 : out std_logic;
    FO157 : out std_logic;
    FO158 : out std_logic;
    FO159 : out std_logic;
    FO160 : out std_logic;
    FO161 : out std_logic;
    FO162 : out std_logic;
    FO163 : out std_logic;
    FO164 : out std_logic;
    FO165 : out std_logic;
    FO166 : out std_logic;
    FO167 : out std_logic;
    FO168 : out std_logic;
    FO169 : out std_logic;
    FO170 : out std_logic;
    FO171 : out std_logic;
    FO172 : out std_logic;
    FO173 : out std_logic;
    FO174 : out std_logic;
    FO175 : out std_logic;
    FO176 : out std_logic;
    FO177 : out std_logic;
    FO178 : out std_logic;
    FO179 : out std_logic;
    FO180 : out std_logic;
    FO181 : out std_logic;
    FO182 : out std_logic;
    FO183 : out std_logic;
    FO184 : out std_logic;
    FO185 : out std_logic;
    FO186 : out std_logic;
    FO187 : out std_logic;
    FO188 : out std_logic;
    FO189 : out std_logic;
    FO190 : out std_logic;
    FO191 : out std_logic;
    FO192 : out std_logic
);
end component NX_RB;

begin

rb: NX_RB
generic map (
    inputClk      => inputClk,
    inputBypass   => inputBypass,
    inputContext  => inputContext,
    outputClk     => outputClk,
    outputBypass  => outputBypass,
    outputContext => outputContext
)
port map (
    CK1   => CK(0),
    CK2   => CK(1),
    CK3   => CK(2),
    CK4   => CK(3),
    EI1   => EI(0),
    EI2   => EI(1),
    EI3   => EI(2),
    EI4   => EI(3),
    EI5   => EI(4),
    EI6   => EI(5),
    EI7   => EI(6),
    EI8   => EI(7),
    EI9   => EI(8),
    EI10  => EI(9),
    EI11  => EI(10),
    EI12  => EI(11),
    EI13  => EI(12),
    EI14  => EI(13),
    EI15  => EI(14),
    EI16  => EI(15),
    EI17  => EI(16),
    EI18  => EI(17),
    EI19  => EI(18),
    EI20  => EI(19),
    EI21  => EI(20),
    EI22  => EI(21),
    EI23  => EI(22),
    EI24  => EI(23),
    EI25  => EI(24),
    EI26  => EI(25),
    EI27  => EI(26),
    EI28  => EI(27),
    EI29  => EI(28),
    EI30  => EI(29),
    EI31  => EI(30),
    EI32  => EI(31),
    EI33  => EI(32),
    EI34  => EI(33),
    EI35  => EI(34),
    EI36  => EI(35),
    EI37  => EI(36),
    EI38  => EI(37),
    EI39  => EI(38),
    EI40  => EI(39),
    EI41  => EI(40),
    EI42  => EI(41),
    EI43  => EI(42),
    EI44  => EI(43),
    EI45  => EI(44),
    EI46  => EI(45),
    EI47  => EI(46),
    EI48  => EI(47),
    EI49  => EI(48),
    EI50  => EI(49),
    EI51  => EI(50),
    EI52  => EI(51),
    EI53  => EI(52),
    EI54  => EI(53),
    EI55  => EI(54),
    EI56  => EI(55),
    EI57  => EI(56),
    EI58  => EI(57),
    EI59  => EI(58),
    EI60  => EI(59),
    EI61  => EI(60),
    EI62  => EI(61),
    EI63  => EI(62),
    EI64  => EI(63),
    EI65  => EI(64),
    EI66  => EI(65),
    EI67  => EI(66),
    EI68  => EI(67),
    EI69  => EI(68),
    EI70  => EI(69),
    EI71  => EI(70),
    EI72  => EI(71),
    EI73  => EI(72),
    EI74  => EI(73),
    EI75  => EI(74),
    EI76  => EI(75),
    EI77  => EI(76),
    EI78  => EI(77),
    EI79  => EI(78),
    EI80  => EI(79),
    EI81  => EI(80),
    EI82  => EI(81),
    EI83  => EI(82),
    EI84  => EI(83),
    EI85  => EI(84),
    EI86  => EI(85),
    EI87  => EI(86),
    EI88  => EI(87),
    EI89  => EI(88),
    EI90  => EI(89),
    EI91  => EI(90),
    EI92  => EI(91),
    EI93  => EI(92),
    EI94  => EI(93),
    EI95  => EI(94),
    EI96  => EI(95),
    EI97  => EI(96),
    EI98  => EI(97),
    EI99  => EI(98),
    EI100 => EI(99),
    EI101 => EI(100),
    EI102 => EI(101),
    EI103 => EI(102),
    EI104 => EI(103),
    EI105 => EI(104),
    EI106 => EI(105),
    EI107 => EI(106),
    EI108 => EI(107),
    EI109 => EI(108),
    EI110 => EI(109),
    EI111 => EI(110),
    EI112 => EI(111),
    EI113 => EI(112),
    EI114 => EI(113),
    EI115 => EI(114),
    EI116 => EI(115),
    EI117 => EI(116),
    EI118 => EI(117),
    EI119 => EI(118),
    EI120 => EI(119),
    EI121 => EI(120),
    EI122 => EI(121),
    EI123 => EI(122),
    EI124 => EI(123),
    EI125 => EI(124),
    EI126 => EI(125),
    EI127 => EI(126),
    EI128 => EI(127),
    EI129 => EI(128),
    EI130 => EI(129),
    EI131 => EI(130),
    EI132 => EI(131),
    EI133 => EI(132),
    EI134 => EI(133),
    EI135 => EI(134),
    EI136 => EI(135),
    EI137 => EI(136),
    EI138 => EI(137),
    EI139 => EI(138),
    EI140 => EI(139),
    EI141 => EI(140),
    EI142 => EI(141),
    EI143 => EI(142),
    EI144 => EI(143),
    EI145 => EI(144),
    EI146 => EI(145),
    EI147 => EI(146),
    EI148 => EI(147),
    EI149 => EI(148),
    EI150 => EI(149),
    EI151 => EI(150),
    EI152 => EI(151),
    EI153 => EI(152),
    EI154 => EI(153),
    EI155 => EI(154),
    EI156 => EI(155),
    EI157 => EI(156),
    EI158 => EI(157),
    EI159 => EI(158),
    EI160 => EI(159),
    EI161 => EI(160),
    EI162 => EI(161),
    EI163 => EI(162),
    EI164 => EI(163),
    EI165 => EI(164),
    EI166 => EI(165),
    EI167 => EI(166),
    EI168 => EI(167),
    EI169 => EI(168),
    EI170 => EI(169),
    EI171 => EI(170),
    EI172 => EI(171),
    EI173 => EI(172),
    EI174 => EI(173),
    EI175 => EI(174),
    EI176 => EI(175),
    EI177 => EI(176),
    EI178 => EI(177),
    EI179 => EI(178),
    EI180 => EI(179),
    EI181 => EI(180),
    EI182 => EI(181),
    EI183 => EI(182),
    EI184 => EI(183),
    EI185 => EI(184),
    EI186 => EI(185),
    EI187 => EI(186),
    EI188 => EI(187),
    EI189 => EI(188),
    EI190 => EI(189),
    EI191 => EI(190),
    EI192 => EI(191),
    EI_CK => EI_CK,
    EO_CK => EO_CK,
    EO1   => EO(0),
    EO2   => EO(1),
    EO3   => EO(2),
    EO4   => EO(3),
    EO5   => EO(4),
    EO6   => EO(5),
    EO7   => EO(6),
    EO8   => EO(7),
    EO9   => EO(8),
    EO10  => EO(9),
    EO11  => EO(10),
    EO12  => EO(11),
    EO13  => EO(12),
    EO14  => EO(13),
    EO15  => EO(14),
    EO16  => EO(15),
    EO17  => EO(16),
    EO18  => EO(17),
    EO19  => EO(18),
    EO20  => EO(19),
    EO21  => EO(20),
    EO22  => EO(21),
    EO23  => EO(22),
    EO24  => EO(23),
    EO25  => EO(24),
    EO26  => EO(25),
    EO27  => EO(26),
    EO28  => EO(27),
    EO29  => EO(28),
    EO30  => EO(29),
    EO31  => EO(30),
    EO32  => EO(31),
    EO33  => EO(32),
    EO34  => EO(33),
    EO35  => EO(34),
    EO36  => EO(35),
    EO37  => EO(36),
    EO38  => EO(37),
    EO39  => EO(38),
    EO40  => EO(39),
    EO41  => EO(40),
    EO42  => EO(41),
    EO43  => EO(42),
    EO44  => EO(43),
    EO45  => EO(44),
    EO46  => EO(45),
    EO47  => EO(46),
    EO48  => EO(47),
    EO49  => EO(48),
    EO50  => EO(49),
    EO51  => EO(50),
    EO52  => EO(51),
    EO53  => EO(52),
    EO54  => EO(53),
    EO55  => EO(54),
    EO56  => EO(55),
    EO57  => EO(56),
    EO58  => EO(57),
    EO59  => EO(58),
    EO60  => EO(59),
    EO61  => EO(60),
    EO62  => EO(61),
    EO63  => EO(62),
    EO64  => EO(63),
    EO65  => EO(64),
    EO66  => EO(65),
    EO67  => EO(66),
    EO68  => EO(67),
    EO69  => EO(68),
    EO70  => EO(69),
    EO71  => EO(70),
    EO72  => EO(71),
    EO73  => EO(72),
    EO74  => EO(73),
    EO75  => EO(74),
    EO76  => EO(75),
    EO77  => EO(76),
    EO78  => EO(77),
    EO79  => EO(78),
    EO80  => EO(79),
    EO81  => EO(80),
    EO82  => EO(81),
    EO83  => EO(82),
    EO84  => EO(83),
    EO85  => EO(84),
    EO86  => EO(85),
    EO87  => EO(86),
    EO88  => EO(87),
    EO89  => EO(88),
    EO90  => EO(89),
    EO91  => EO(90),
    EO92  => EO(91),
    EO93  => EO(92),
    EO94  => EO(93),
    EO95  => EO(94),
    EO96  => EO(95),
    EO97  => EO(96),
    EO98  => EO(97),
    EO99  => EO(98),
    EO100 => EO(99),
    EO101 => EO(100),
    EO102 => EO(101),
    EO103 => EO(102),
    EO104 => EO(103),
    EO105 => EO(104),
    EO106 => EO(105),
    EO107 => EO(106),
    EO108 => EO(107),
    EO109 => EO(108),
    EO110 => EO(109),
    EO111 => EO(110),
    EO112 => EO(111),
    EO113 => EO(112),
    EO114 => EO(113),
    EO115 => EO(114),
    EO116 => EO(115),
    EO117 => EO(116),
    EO118 => EO(117),
    EO119 => EO(118),
    EO120 => EO(119),
    EO121 => EO(120),
    EO122 => EO(121),
    EO123 => EO(122),
    EO124 => EO(123),
    EO125 => EO(124),
    EO126 => EO(125),
    EO127 => EO(126),
    EO128 => EO(127),
    EO129 => EO(128),
    EO130 => EO(129),
    EO131 => EO(130),
    EO132 => EO(131),
    EO133 => EO(132),
    EO134 => EO(133),
    EO135 => EO(134),
    EO136 => EO(135),
    EO137 => EO(136),
    EO138 => EO(137),
    EO139 => EO(138),
    EO140 => EO(139),
    EO141 => EO(140),
    EO142 => EO(141),
    EO143 => EO(142),
    EO144 => EO(143),
    EO145 => EO(144),
    EO146 => EO(145),
    EO147 => EO(146),
    EO148 => EO(147),
    EO149 => EO(148),
    EO150 => EO(149),
    EO151 => EO(150),
    EO152 => EO(151),
    EO153 => EO(152),
    EO154 => EO(153),
    EO155 => EO(154),
    EO156 => EO(155),
    EO157 => EO(156),
    EO158 => EO(157),
    EO159 => EO(158),
    EO160 => EO(159),
    EO161 => EO(160),
    EO162 => EO(161),
    EO163 => EO(162),
    EO164 => EO(163),
    EO165 => EO(164),
    EO166 => EO(165),
    EO167 => EO(166),
    EO168 => EO(167),
    EO169 => EO(168),
    EO170 => EO(169),
    EO171 => EO(170),
    EO172 => EO(171),
    EO173 => EO(172),
    EO174 => EO(173),
    EO175 => EO(174),
    EO176 => EO(175),
    EO177 => EO(176),
    EO178 => EO(177),
    EO179 => EO(178),
    EO180 => EO(179),
    EO181 => EO(180),
    EO182 => EO(181),
    EO183 => EO(182),
    EO184 => EO(183),
    EO185 => EO(184),
    EO186 => EO(185),
    EO187 => EO(186),
    EO188 => EO(187),
    EO189 => EO(188),
    EO190 => EO(189),
    EO191 => EO(190),
    EO192 => EO(191),
    FI1   => FI(0),
    FI2   => FI(1),
    FI3   => FI(2),
    FI4   => FI(3),
    FI5   => FI(4),
    FI6   => FI(5),
    FI7   => FI(6),
    FI8   => FI(7),
    FI9   => FI(8),
    FI10  => FI(9),
    FI11  => FI(10),
    FI12  => FI(11),
    FI13  => FI(12),
    FI14  => FI(13),
    FI15  => FI(14),
    FI16  => FI(15),
    FI17  => FI(16),
    FI18  => FI(17),
    FI19  => FI(18),
    FI20  => FI(19),
    FI21  => FI(20),
    FI22  => FI(21),
    FI23  => FI(22),
    FI24  => FI(23),
    FI25  => FI(24),
    FI26  => FI(25),
    FI27  => FI(26),
    FI28  => FI(27),
    FI29  => FI(28),
    FI30  => FI(29),
    FI31  => FI(30),
    FI32  => FI(31),
    FI33  => FI(32),
    FI34  => FI(33),
    FI35  => FI(34),
    FI36  => FI(35),
    FI37  => FI(36),
    FI38  => FI(37),
    FI39  => FI(38),
    FI40  => FI(39),
    FI41  => FI(40),
    FI42  => FI(41),
    FI43  => FI(42),
    FI44  => FI(43),
    FI45  => FI(44),
    FI46  => FI(45),
    FI47  => FI(46),
    FI48  => FI(47),
    FI49  => FI(48),
    FI50  => FI(49),
    FI51  => FI(50),
    FI52  => FI(51),
    FI53  => FI(52),
    FI54  => FI(53),
    FI55  => FI(54),
    FI56  => FI(55),
    FI57  => FI(56),
    FI58  => FI(57),
    FI59  => FI(58),
    FI60  => FI(59),
    FI61  => FI(60),
    FI62  => FI(61),
    FI63  => FI(62),
    FI64  => FI(63),
    FI65  => FI(64),
    FI66  => FI(65),
    FI67  => FI(66),
    FI68  => FI(67),
    FI69  => FI(68),
    FI70  => FI(69),
    FI71  => FI(70),
    FI72  => FI(71),
    FI73  => FI(72),
    FI74  => FI(73),
    FI75  => FI(74),
    FI76  => FI(75),
    FI77  => FI(76),
    FI78  => FI(77),
    FI79  => FI(78),
    FI80  => FI(79),
    FI81  => FI(80),
    FI82  => FI(81),
    FI83  => FI(82),
    FI84  => FI(83),
    FI85  => FI(84),
    FI86  => FI(85),
    FI87  => FI(86),
    FI88  => FI(87),
    FI89  => FI(88),
    FI90  => FI(89),
    FI91  => FI(90),
    FI92  => FI(91),
    FI93  => FI(92),
    FI94  => FI(93),
    FI95  => FI(94),
    FI96  => FI(95),
    FI97  => FI(96),
    FI98  => FI(97),
    FI99  => FI(98),
    FI100 => FI(99),
    FI101 => FI(100),
    FI102 => FI(101),
    FI103 => FI(102),
    FI104 => FI(103),
    FI105 => FI(104),
    FI106 => FI(105),
    FI107 => FI(106),
    FI108 => FI(107),
    FI109 => FI(108),
    FI110 => FI(109),
    FI111 => FI(110),
    FI112 => FI(111),
    FI113 => FI(112),
    FI114 => FI(113),
    FI115 => FI(114),
    FI116 => FI(115),
    FI117 => FI(116),
    FI118 => FI(117),
    FI119 => FI(118),
    FI120 => FI(119),
    FI121 => FI(120),
    FI122 => FI(121),
    FI123 => FI(122),
    FI124 => FI(123),
    FI125 => FI(124),
    FI126 => FI(125),
    FI127 => FI(126),
    FI128 => FI(127),
    FI129 => FI(128),
    FI130 => FI(129),
    FI131 => FI(130),
    FI132 => FI(131),
    FI133 => FI(132),
    FI134 => FI(133),
    FI135 => FI(134),
    FI136 => FI(135),
    FI137 => FI(136),
    FI138 => FI(137),
    FI139 => FI(138),
    FI140 => FI(139),
    FI141 => FI(140),
    FI142 => FI(141),
    FI143 => FI(142),
    FI144 => FI(143),
    FI145 => FI(144),
    FI146 => FI(145),
    FI147 => FI(146),
    FI148 => FI(147),
    FI149 => FI(148),
    FI150 => FI(149),
    FI151 => FI(150),
    FI152 => FI(151),
    FI153 => FI(152),
    FI154 => FI(153),
    FI155 => FI(154),
    FI156 => FI(155),
    FI157 => FI(156),
    FI158 => FI(157),
    FI159 => FI(158),
    FI160 => FI(159),
    FI161 => FI(160),
    FI162 => FI(161),
    FI163 => FI(162),
    FI164 => FI(163),
    FI165 => FI(164),
    FI166 => FI(165),
    FI167 => FI(166),
    FI168 => FI(167),
    FI169 => FI(168),
    FI170 => FI(169),
    FI171 => FI(170),
    FI172 => FI(171),
    FI173 => FI(172),
    FI174 => FI(173),
    FI175 => FI(174),
    FI176 => FI(175),
    FI177 => FI(176),
    FI178 => FI(177),
    FI179 => FI(178),
    FI180 => FI(179),
    FI181 => FI(180),
    FI182 => FI(181),
    FI183 => FI(182),
    FI184 => FI(183),
    FI185 => FI(184),
    FI186 => FI(185),
    FI187 => FI(186),
    FI188 => FI(187),
    FI189 => FI(188),
    FI190 => FI(189),
    FI191 => FI(190),
    FI192 => FI(191),
    FO1   => FO(0),
    FO2   => FO(1),
    FO3   => FO(2),
    FO4   => FO(3),
    FO5   => FO(4),
    FO6   => FO(5),
    FO7   => FO(6),
    FO8   => FO(7),
    FO9   => FO(8),
    FO10  => FO(9),
    FO11  => FO(10),
    FO12  => FO(11),
    FO13  => FO(12),
    FO14  => FO(13),
    FO15  => FO(14),
    FO16  => FO(15),
    FO17  => FO(16),
    FO18  => FO(17),
    FO19  => FO(18),
    FO20  => FO(19),
    FO21  => FO(20),
    FO22  => FO(21),
    FO23  => FO(22),
    FO24  => FO(23),
    FO25  => FO(24),
    FO26  => FO(25),
    FO27  => FO(26),
    FO28  => FO(27),
    FO29  => FO(28),
    FO30  => FO(29),
    FO31  => FO(30),
    FO32  => FO(31),
    FO33  => FO(32),
    FO34  => FO(33),
    FO35  => FO(34),
    FO36  => FO(35),
    FO37  => FO(36),
    FO38  => FO(37),
    FO39  => FO(38),
    FO40  => FO(39),
    FO41  => FO(40),
    FO42  => FO(41),
    FO43  => FO(42),
    FO44  => FO(43),
    FO45  => FO(44),
    FO46  => FO(45),
    FO47  => FO(46),
    FO48  => FO(47),
    FO49  => FO(48),
    FO50  => FO(49),
    FO51  => FO(50),
    FO52  => FO(51),
    FO53  => FO(52),
    FO54  => FO(53),
    FO55  => FO(54),
    FO56  => FO(55),
    FO57  => FO(56),
    FO58  => FO(57),
    FO59  => FO(58),
    FO60  => FO(59),
    FO61  => FO(60),
    FO62  => FO(61),
    FO63  => FO(62),
    FO64  => FO(63),
    FO65  => FO(64),
    FO66  => FO(65),
    FO67  => FO(66),
    FO68  => FO(67),
    FO69  => FO(68),
    FO70  => FO(69),
    FO71  => FO(70),
    FO72  => FO(71),
    FO73  => FO(72),
    FO74  => FO(73),
    FO75  => FO(74),
    FO76  => FO(75),
    FO77  => FO(76),
    FO78  => FO(77),
    FO79  => FO(78),
    FO80  => FO(79),
    FO81  => FO(80),
    FO82  => FO(81),
    FO83  => FO(82),
    FO84  => FO(83),
    FO85  => FO(84),
    FO86  => FO(85),
    FO87  => FO(86),
    FO88  => FO(87),
    FO89  => FO(88),
    FO90  => FO(89),
    FO91  => FO(90),
    FO92  => FO(91),
    FO93  => FO(92),
    FO94  => FO(93),
    FO95  => FO(94),
    FO96  => FO(95),
    FO97  => FO(96),
    FO98  => FO(97),
    FO99  => FO(98),
    FO100 => FO(99),
    FO101 => FO(100),
    FO102 => FO(101),
    FO103 => FO(102),
    FO104 => FO(103),
    FO105 => FO(104),
    FO106 => FO(105),
    FO107 => FO(106),
    FO108 => FO(107),
    FO109 => FO(108),
    FO110 => FO(109),
    FO111 => FO(110),
    FO112 => FO(111),
    FO113 => FO(112),
    FO114 => FO(113),
    FO115 => FO(114),
    FO116 => FO(115),
    FO117 => FO(116),
    FO118 => FO(117),
    FO119 => FO(118),
    FO120 => FO(119),
    FO121 => FO(120),
    FO122 => FO(121),
    FO123 => FO(122),
    FO124 => FO(123),
    FO125 => FO(124),
    FO126 => FO(125),
    FO127 => FO(126),
    FO128 => FO(127),
    FO129 => FO(128),
    FO130 => FO(129),
    FO131 => FO(130),
    FO132 => FO(131),
    FO133 => FO(132),
    FO134 => FO(133),
    FO135 => FO(134),
    FO136 => FO(135),
    FO137 => FO(136),
    FO138 => FO(137),
    FO139 => FO(138),
    FO140 => FO(139),
    FO141 => FO(140),
    FO142 => FO(141),
    FO143 => FO(142),
    FO144 => FO(143),
    FO145 => FO(144),
    FO146 => FO(145),
    FO147 => FO(146),
    FO148 => FO(147),
    FO149 => FO(148),
    FO150 => FO(149),
    FO151 => FO(150),
    FO152 => FO(151),
    FO153 => FO(152),
    FO154 => FO(153),
    FO155 => FO(154),
    FO156 => FO(155),
    FO157 => FO(156),
    FO158 => FO(157),
    FO159 => FO(158),
    FO160 => FO(159),
    FO161 => FO(160),
    FO162 => FO(161),
    FO163 => FO(162),
    FO164 => FO(163),
    FO165 => FO(164),
    FO166 => FO(165),
    FO167 => FO(166),
    FO168 => FO(167),
    FO169 => FO(168),
    FO170 => FO(169),
    FO171 => FO(170),
    FO172 => FO(171),
    FO173 => FO(172),
    FO174 => FO(173),
    FO175 => FO(174),
    FO176 => FO(175),
    FO177 => FO(176),
    FO178 => FO(177),
    FO179 => FO(178),
    FO180 => FO(179),
    FO181 => FO(180),
    FO182 => FO(181),
    FO183 => FO(182),
    FO184 => FO(183),
    FO185 => FO(184),
    FO186 => FO(185),
    FO187 => FO(186),
    FO188 => FO(187),
    FO189 => FO(188),
    FO190 => FO(189),
    FO191 => FO(190),
    FO192 => FO(191)
);
end NX_RTL;

-- =================================================================================================
--   NX_RFB_L definition                                                                2017/09/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_RFB_L is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic;
    XRCK : out std_logic;
    XRO1 : out std_logic;
    XRO2 : out std_logic;
    XRO3 : out std_logic;
    XRO4 : out std_logic;
    XRO5 : out std_logic;
    XRO6 : out std_logic;
    XWCK : out std_logic;
    XWO1 : out std_logic;
    XWO2 : out std_logic;
    XWO3 : out std_logic;
    XWO4 : out std_logic;
    XWO5 : out std_logic;
    XWO6 : out std_logic
);
end NX_RFB_L;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RFB_L_WRAP definition                                                           2017/09/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_RFB_L_WRAP is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I   : in  std_logic_vector(15 downto 0);
    COR : out std_logic;
    ERR : out std_logic;
    O   : out std_logic_vector(15 downto 0);
    RA  : in  std_logic_vector(5 downto 0);
    RE  : in  std_logic;
    WA  : in  std_logic_vector(5 downto 0);
    WE  : in  std_logic;
    XRCK : out std_logic;
    XRO  : out std_logic_vector(5 downto 0);
    XWCK : out std_logic;
    XWO  : out std_logic_vector(5 downto 0)
);
end NX_RFB_L_WRAP;

architecture NX_RTL of NX_RFB_L_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_L
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic;
    XRCK : out std_logic;
    XRO1 : out std_logic;
    XRO2 : out std_logic;
    XRO3 : out std_logic;
    XRO4 : out std_logic;
    XRO5 : out std_logic;
    XRO6 : out std_logic;
    XWCK : out std_logic;
    XWO1 : out std_logic;
    XWO2 : out std_logic;
    XWO3 : out std_logic;
    XWO4 : out std_logic;
    XWO5 : out std_logic;
    XWO6 : out std_logic
);
end component NX_RFB_L;

begin

rfb: NX_RFB_L generic map (
    rck_edge    => rck_edge,
    wck_edge    => wck_edge,
    mem_ctxt    => mem_ctxt)
port map (
    RCK => RCK,
    WCK => WCK,
    I1  => I(0),
    I2  => I(1),
    I3  => I(2),
    I4  => I(3),
    I5  => I(4),
    I6  => I(5),
    I7  => I(6),
    I8  => I(7),
    I9  => I(8),
    I10 => I(9),
    I11 => I(10),
    I12 => I(11),
    I13 => I(12),
    I14 => I(13),
    I15 => I(14),
    I16 => I(15),
    COR => COR,
    ERR => ERR,
    O1  => O(0),
    O2  => O(1),
    O3  => O(2),
    O4  => O(3),
    O5  => O(4),
    O6  => O(5),
    O7  => O(6),
    O8  => O(7),
    O9  => O(8),
    O10 => O(9),
    O11 => O(10),
    O12 => O(11),
    O13 => O(12),
    O14 => O(13),
    O15 => O(14),
    O16 => O(15),
    RA1 => RA(0),
    RA2 => RA(1),
    RA3 => RA(2),
    RA4 => RA(3),
    RA5 => RA(4),
    RA6 => RA(5),
    RE  => RE,
    WA1 => WA(0),
    WA2 => WA(1),
    WA3 => WA(2),
    WA4 => WA(3),
    WA5 => WA(4),
    WA6 => WA(5),
    WE  => WE,
    XRCK => XRCK,
    XRO1 => XRO(0),
    XRO2 => XRO(1),
    XRO3 => XRO(2),
    XRO4 => XRO(3),
    XRO5 => XRO(4),
    XRO6 => XRO(5),
    XWCK => XWCK,
    XWO1 => XWO(0),
    XWO2 => XWO(1),
    XWO3 => XWO(2),
    XWO4 => XWO(3),
    XWO5 => XWO(4),
    XWO6 => XWO(5)
);
end NX_RTL;
-- =================================================================================================
--   NX_RFB_M definition                                                                 2017/09/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_RFB_M is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic
);
end NX_RFB_M;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RFB_WRAP definition                                                             2017/09/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_RFB_WRAP is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I   : in  std_logic_vector(15 downto 0);
    COR : out std_logic;
    ERR : out std_logic;
    O   : out std_logic_vector(15 downto 0);
    RA  : in  std_logic_vector(5 downto 0);
    RE  : in  std_logic;
    WA  : in  std_logic_vector(5 downto 0);
    WE  : in  std_logic
);
end NX_RFB_WRAP;

architecture NX_RTL of NX_RFB_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_M
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic
);
end component NX_RFB_M;

begin

rfb: NX_RFB_M generic map (
    rck_edge    => rck_edge,
    wck_edge    => wck_edge,
    mem_ctxt    => mem_ctxt)
port map (
    RCK => RCK,
    WCK => WCK,
    I1  => I(0),
    I2  => I(1),
    I3  => I(2),
    I4  => I(3),
    I5  => I(4),
    I6  => I(5),
    I7  => I(6),
    I8  => I(7),
    I9  => I(8),
    I10 => I(9),
    I11 => I(10),
    I12 => I(11),
    I13 => I(12),
    I14 => I(13),
    I15 => I(14),
    I16 => I(15),
    COR => COR,
    ERR => ERR,
    O1  => O(0),
    O2  => O(1),
    O3  => O(2),
    O4  => O(3),
    O5  => O(4),
    O6  => O(5),
    O7  => O(6),
    O8  => O(7),
    O9  => O(8),
    O10 => O(9),
    O11 => O(10),
    O12 => O(11),
    O13 => O(12),
    O14 => O(13),
    O15 => O(14),
    O16 => O(15),
    RA1 => RA(0),
    RA2 => RA(1),
    RA3 => RA(2),
    RA4 => RA(3),
    RA5 => RA(4),
    RA6 => RA(5),
    RE  => RE,
    WA1 => WA(0),
    WA2 => WA(1),
    WA3 => WA(2),
    WA4 => WA(3),
    WA5 => WA(4),
    WA6 => WA(5),
    WE  => WE
);
end NX_RTL;

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_CKS is
port (
    CKI : in  std_logic;
    CMD : in  std_logic;
    CKO : out std_logic
);
end NX_CKS;
-- =================================================================================================
--   NX_RFB (compatible) definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_RFB is
generic (
    rck_edge  : bit := '0';   -- 0: read  clock rising edge - 1: read  clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic
);
end NX_RFB;

architecture NX_RTL of NX_RFB is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_M is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic
);
end component NX_RFB_M;

component NX_RFB_L is
generic (
    rck_edge  : bit := '0';   -- 0: read clock rising edge - 1: read clock falling edge
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    RCK : in  std_logic;
    WCK : in  std_logic;
    I1  : in  std_logic;
    I2  : in  std_logic;
    I3  : in  std_logic;
    I4  : in  std_logic;
    I5  : in  std_logic;
    I6  : in  std_logic;
    I7  : in  std_logic;
    I8  : in  std_logic;
    I9  : in  std_logic;
    I10 : in  std_logic;
    I11 : in  std_logic;
    I12 : in  std_logic;
    I13 : in  std_logic;
    I14 : in  std_logic;
    I15 : in  std_logic;
    I16 : in  std_logic;
    COR : out std_logic;
    ERR : out std_logic;
    O1  : out std_logic;
    O2  : out std_logic;
    O3  : out std_logic;
    O4  : out std_logic;
    O5  : out std_logic;
    O6  : out std_logic;
    O7  : out std_logic;
    O8  : out std_logic;
    O9  : out std_logic;
    O10 : out std_logic;
    O11 : out std_logic;
    O12 : out std_logic;
    O13 : out std_logic;
    O14 : out std_logic;
    O15 : out std_logic;
    O16 : out std_logic;
    RA1 : in  std_logic;
    RA2 : in  std_logic;
    RA3 : in  std_logic;
    RA4 : in  std_logic;
    RA5 : in  std_logic;
    RA6 : in  std_logic;
    RE  : in  std_logic;
    WA1 : in  std_logic;
    WA2 : in  std_logic;
    WA3 : in  std_logic;
    WA4 : in  std_logic;
    WA5 : in  std_logic;
    WA6 : in  std_logic;
    WE  : in  std_logic;
    XRCK : out std_logic;
    XRO1 : out std_logic;
    XRO2 : out std_logic;
    XRO3 : out std_logic;
    XRO4 : out std_logic;
    XRO5 : out std_logic;
    XRO6 : out std_logic;
    XWCK : out std_logic;
    XWO1 : out std_logic;
    XWO2 : out std_logic;
    XWO3 : out std_logic;
    XWO4 : out std_logic;
    XWO5 : out std_logic;
    XWO6 : out std_logic
);
end component NX_RFB_L;

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

component NX_DFF is
generic (
    dff_edge   : bit := '0';
    dff_init   : bit := '0';
    dff_load   : bit := '0';
    dff_sync   : bit := '0';
    dff_ctxt   : std_logic := 'U'
);
port (
    I  : in  std_logic;
    CK : in  std_logic;
    L  : in  std_logic;
    R  : in  std_logic;
    O  : out std_logic
);
end component NX_DFF;

begin

medium : if NX_SYMBOL = "NG_M" generate
    rfb: NX_RFB_M generic map (
        rck_edge    => rck_edge,
        wck_edge    => wck_edge,
        mem_ctxt    => mem_ctxt)
    port map (
        RCK => RCK,
        WCK => WCK,
        I1  => I1,
        I2  => I2,
        I3  => I3,
        I4  => I4,
        I5  => I5,
        I6  => I6,
        I7  => I7,
        I8  => I8,
        I9  => I9,
        I10 => I10,
        I11 => I11,
        I12 => I12,
        I13 => I13,
        I14 => I14,
        I15 => I15,
        I16 => I16,
        COR => COR,
        ERR => ERR,
        O1  => O1,
        O2  => O2,
        O3  => O3,
        O4  => O4,
        O5  => O5,
        O6  => O6,
        O7  => O7,
        O8  => O8,
        O9  => O9,
        O10 => O10,
        O11 => O11,
        O12 => O12,
        O13 => O13,
        O14 => O14,
        O15 => O15,
        O16 => O16,
        RA1 => RA1,
        RA2 => RA2,
        RA3 => RA3,
        RA4 => RA4,
        RA5 => RA5,
        RA6 => RA6,
        RE  => RE,
        WA1 => WA1,
        WA2 => WA2,
        WA3 => WA3,
        WA4 => WA4,
        WA5 => WA5,
        WA6 => WA6,
        WE  => WE
    );
end generate;

large : if NX_SYMBOL = "NG_L" generate
    rfb: NX_RFB_L generic map (
        rck_edge    => rck_edge,
        wck_edge    => wck_edge,
        mem_ctxt    => mem_ctxt)
    port map (
        RCK => RCK,
        WCK => WCK,
        I1  => I1,
        I2  => I2,
        I3  => I3,
        I4  => I4,
        I5  => I5,
        I6  => I6,
        I7  => I7,
        I8  => I8,
        I9  => I9,
        I10 => I10,
        I11 => I11,
        I12 => I12,
        I13 => I13,
        I14 => I14,
        I15 => I15,
        I16 => I16,
        COR => COR,
        ERR => ERR,
        O1  => O1,
        O2  => O2,
        O3  => O3,
        O4  => O4,
        O5  => O5,
        O6  => O6,
        O7  => O7,
        O8  => O8,
        O9  => O9,
        O10 => O10,
        O11 => O11,
        O12 => O12,
        O13 => O13,
        O14 => O14,
        O15 => O15,
        O16 => O16,
        RA1 => RA1,
        RA2 => RA2,
        RA3 => RA3,
        RA4 => RA4,
        RA5 => RA5,
        RA6 => RA6,
        RE  => RE,
        WA1 => WA1,
        WA2 => WA2,
        WA3 => WA3,
        WA4 => WA4,
        WA5 => WA5,
        WA6 => WA6,
        WE  => WE,
        XRCK => OPEN,
        XRO1 => OPEN,
        XRO2 => OPEN,
        XRO3 => OPEN,
        XRO4 => OPEN,
        XRO5 => OPEN,
        XRO6 => OPEN,
        XWCK => OPEN,
        XWO1 => OPEN,
        XWO2 => OPEN,
        XWO3 => OPEN,
        XWO4 => OPEN,
        XWO5 => OPEN,
        XWO6 => OPEN
    );
end generate;

ultra : if NX_SYMBOL = "NG_U" or NX_SYMBOL = "NG_C" generate
signal D : std_logic_vector(15 downto 0);
signal Q : std_logic_vector(15 downto 0);

begin
rfb: NX_RFB_U
generic map (
    mode      => 2, -- 2: DPREG_64x18
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I1,
    I2   => I2,
    I3   => I3,
    I4   => I4,
    I5   => I5,
    I6   => I6,
    I7   => I7,
    I8   => I8,
    I9   => I9,
    I10  => I10,
    I11  => I11,
    I12  => I12,
    I13  => I13,
    I14  => I14,
    I15  => I15,
    I16  => I16,
    I17  => '0',
    I18  => '0',
    I19  => '0',
    I20  => '0',
    I21  => '0',
    I22  => '0',
    I23  => '0',
    I24  => '0',
    I25  => '0',
    I26  => '0',
    I27  => '0',
    I28  => '0',
    I29  => '0',
    I30  => '0',
    I31  => '0',
    I32  => '0',
    I33  => '0',
    I34  => '0',
    I35  => '0',
    I36  => '0',
    O1   => D(0),
    O2   => D(1),
    O3   => D(2),
    O4   => D(3),
    O5   => D(4),
    O6   => D(5),
    O7   => D(6),
    O8   => D(7),
    O9   => D(8),
    O10  => D(9),
    O11  => D(10),
    O12  => D(11),
    O13  => D(12),
    O14  => D(13),
    O15  => D(14),
    O16  => D(15),
    O17  => OPEN,
    O18  => OPEN,
    O19  => OPEN,
    O20  => OPEN,
    O21  => OPEN,
    O22  => OPEN,
    O23  => OPEN,
    O24  => OPEN,
    O25  => OPEN,
    O26  => OPEN,
    O27  => OPEN,
    O28  => OPEN,
    O29  => OPEN,
    O30  => OPEN,
    O31  => OPEN,
    O32  => OPEN,
    O33  => OPEN,
    O34  => OPEN,
    O35  => OPEN,
    O36  => OPEN,
    RA1  => RA1,
    RA2  => RA2,
    RA3  => RA3,
    RA4  => RA4,
    RA5  => RA5,
    RA6  => RA6,
    RA7  => '0',
    RA8  => '0',
    RA9  => '0',
    RA10 => '0',
    WA1  => WA1,
    WA2  => WA2,
    WA3  => WA3,
    WA4  => WA4,
    WA5  => WA5,
    WA6  => WA6,
    WE   => WE,
    WEA  => '0'
);

OUT_REG : for I in Q'range generate

    reg : NX_DFF
    generic map (
	dff_edge => rck_edge,
	dff_init => '0',
	dff_load => '1'
    )
    port map (
	CK => RCK,
	I  => D(I),
	L  => RE,
	R  => '0',
	O  => Q(I)
    );

end generate;

O1   <= Q(0);
O2   <= Q(1);
O3   <= Q(2);
O4   <= Q(3);
O5   <= Q(4);
O6   <= Q(5);
O7   <= Q(6);
O8   <= Q(7);
O9   <= Q(8);
O10  <= Q(9);
O11  <= Q(10);
O12  <= Q(11);
O13  <= Q(12);
O14  <= Q(13);
O15  <= Q(14);
O16  <= Q(15);

COR <= '0';
ERR <= '0';
end generate;
end NX_RTL;
-- =================================================================================================
--   NX_CDC_U_2DFF definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CDC_U_2DFF is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_adest_arst : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ADRSTI : in  std_logic;
    ADRSTO : out std_logic;
    AI     : in  std_logic_vector(5 downto 0);
    AO     : out std_logic_vector(5 downto 0);
    BDRSTI : in  std_logic;
    BDRSTO : out std_logic;
    BI     : in  std_logic_vector(5 downto 0);
    BO     : out std_logic_vector(5 downto 0)
);
end NX_CDC_U_2DFF;

architecture NX_RTL of NX_CDC_U_2DFF is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 0, -- 0: 2DFF
    ck0_edge       => ck0_edge,
    ck1_edge       => ck1_edge,
    ack_sel        => ack_sel,
    bck_sel        => bck_sel,
    cck_sel        => '0',
    dck_sel        => '0',
    use_asrc_arst  => '0',
    use_adest_arst => use_adest_arst,
    use_bsrc_arst  => '0',
    use_bdest_arst => use_bdest_arst,
    use_csrc_arst  => '0',
    use_cdest_arst => '0',
    use_dsrc_arst  => '0',
    use_ddest_arst => '0',
    link_BA        => '0',
    link_CB        => '0',
    link_DC        => '0'
)
port map (
    CK1    => CK1,
    CK2    => CK2,
    ASRSTI => '0',
    ADRSTI => ADRSTI,
    ASRSTO => OPEN,
    ADRSTO => ADRSTO,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => '0',
    BDRSTI => BDRSTI,
    BSRSTO => OPEN,
    BDRSTO => BDRSTO,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => '0',
    CDRSTI => '0',
    CSRSTO => OPEN,
    CDRSTO => OPEN,
    CI1    => '0',
    CI2    => '0',
    CI3    => '0',
    CI4    => '0',
    CI5    => '0',
    CI6    => '0',
    CO1    => OPEN,
    CO2    => OPEN,
    CO3    => OPEN,
    CO4    => OPEN,
    CO5    => OPEN,
    CO6    => OPEN,
    DSRSTI => '0',
    DDRSTI => '0',
    DSRSTO => OPEN,
    DDRSTO => OPEN,
    DI1    => '0',
    DI2    => '0',
    DI3    => '0',
    DI4    => '0',
    DI5    => '0',
    DI6    => '0',
    DO1    => OPEN,
    DO2    => OPEN,
    DO3    => OPEN,
    DO4    => OPEN,
    DO5    => OPEN,
    DO6    => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U_3DFF definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CDC_U_3DFF is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI     : in  std_logic_vector(5 downto 0);
    AO     : out std_logic_vector(5 downto 0);
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI     : in  std_logic_vector(5 downto 0);
    BO     : out std_logic_vector(5 downto 0)
);
end NX_CDC_U_3DFF;

architecture NX_RTL of NX_CDC_U_3DFF is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 1, -- 1: 3DFF
    ck0_edge       => ck0_edge,
    ck1_edge       => ck1_edge,
    ack_sel        => ack_sel,
    bck_sel        => bck_sel,
    cck_sel        => '0',
    dck_sel        => '0',
    use_asrc_arst  => use_asrc_arst,
    use_adest_arst => use_adest_arst,
    use_bsrc_arst  => use_bsrc_arst,
    use_bdest_arst => use_bdest_arst,
    use_csrc_arst  => '0',
    use_cdest_arst => '0',
    use_dsrc_arst  => '0',
    use_ddest_arst => '0',
    link_BA        => '0',
    link_CB        => '0',
    link_DC        => '0'
)
port map (
    CK1    => CK1,
    CK2    => CK2,
    ASRSTI => ASRSTI,
    ADRSTI => ADRSTI,
    ASRSTO => ASRSTO,
    ADRSTO => ADRSTO,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => BSRSTI,
    BDRSTI => BDRSTI,
    BSRSTO => BSRSTO,
    BDRSTO => BDRSTO,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => '0',
    CDRSTI => '0',
    CSRSTO => OPEN,
    CDRSTO => OPEN,
    CI1    => '0',
    CI2    => '0',
    CI3    => '0',
    CI4    => '0',
    CI5    => '0',
    CI6    => '0',
    CO1    => OPEN,
    CO2    => OPEN,
    CO3    => OPEN,
    CO4    => OPEN,
    CO5    => OPEN,
    CO6    => OPEN,
    DSRSTI => '0',
    DDRSTI => '0',
    DSRSTO => OPEN,
    DDRSTO => OPEN,
    DI1    => '0',
    DI2    => '0',
    DI3    => '0',
    DI4    => '0',
    DI5    => '0',
    DI6    => '0',
    DO1    => OPEN,
    DO2    => OPEN,
    DO3    => OPEN,
    DO4    => OPEN,
    DO5    => OPEN,
    DO6    => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U_FULL definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CDC_U_FULL is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI     : in  std_logic_vector(5 downto 0);
    AO     : out std_logic_vector(5 downto 0);
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI     : in  std_logic_vector(5 downto 0);
    BO     : out std_logic_vector(5 downto 0)
);
end NX_CDC_U_FULL;

architecture NX_RTL of NX_CDC_U_FULL is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 2, -- 2: bin2gray + 3DFF + gray2bin
    ck0_edge       => ck0_edge,
    ck1_edge       => ck1_edge,
    ack_sel        => ack_sel,
    bck_sel        => bck_sel,
    cck_sel        => '0',
    dck_sel        => '0',
    use_asrc_arst  => use_asrc_arst,
    use_adest_arst => use_adest_arst,
    use_bsrc_arst  => use_bsrc_arst,
    use_bdest_arst => use_bdest_arst,
    use_csrc_arst  => '0',
    use_cdest_arst => '0',
    use_dsrc_arst  => '0',
    use_ddest_arst => '0',
    link_BA        => '0',
    link_CB        => '0',
    link_DC        => '0'
)
port map (
    CK1    => CK1,
    CK2    => CK2,
    ASRSTI => ASRSTI,
    ADRSTI => ADRSTI,
    ASRSTO => ASRSTO,
    ADRSTO => ADRSTO,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => BSRSTI,
    BDRSTI => BDRSTI,
    BSRSTO => BSRSTO,
    BDRSTO => BDRSTO,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => '0',
    CDRSTI => '0',
    CSRSTO => OPEN,
    CDRSTO => OPEN,
    CI1    => '0',
    CI2    => '0',
    CI3    => '0',
    CI4    => '0',
    CI5    => '0',
    CI6    => '0',
    CO1    => OPEN,
    CO2    => OPEN,
    CO3    => OPEN,
    CO4    => OPEN,
    CO5    => OPEN,
    CO6    => OPEN,
    DSRSTI => '0',
    DDRSTI => '0',
    DSRSTO => OPEN,
    DDRSTO => OPEN,
    DI1    => '0',
    DI2    => '0',
    DI3    => '0',
    DI4    => '0',
    DI5    => '0',
    DI6    => '0',
    DO1    => OPEN,
    DO2    => OPEN,
    DO3    => OPEN,
    DO4    => OPEN,
    DO5    => OPEN,
    DO6    => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U_BIN2GRAY definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CDC_U_BIN2GRAY is
port (
    AI     : in  std_logic_vector(5 downto 0);
    AO     : out std_logic_vector(5 downto 0);
    BI     : in  std_logic_vector(5 downto 0);
    BO     : out std_logic_vector(5 downto 0)
);
end NX_CDC_U_BIN2GRAY;

architecture NX_RTL of NX_CDC_U_BIN2GRAY is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 3, -- 3: bin2gray
    ck0_edge       => '0',
    ck1_edge       => '0',
    ack_sel        => '0',
    bck_sel        => '0',
    cck_sel        => '0',
    dck_sel        => '0',
    use_asrc_arst  => '0',
    use_adest_arst => '0',
    use_bsrc_arst  => '0',
    use_bdest_arst => '0',
    use_csrc_arst  => '0',
    use_cdest_arst => '0',
    use_dsrc_arst  => '0',
    use_ddest_arst => '0',
    link_BA        => '0',
    link_CB        => '0',
    link_DC        => '0'
)
port map (
    CK1    => '0',
    CK2    => '0',
    ASRSTI => '0',
    ADRSTI => '0',
    ASRSTO => OPEN,
    ADRSTO => OPEN,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => '0',
    BDRSTI => '0',
    BSRSTO => OPEN,
    BDRSTO => OPEN,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => '0',
    CDRSTI => '0',
    CSRSTO => OPEN,
    CDRSTO => OPEN,
    CI1    => '0',
    CI2    => '0',
    CI3    => '0',
    CI4    => '0',
    CI5    => '0',
    CI6    => '0',
    CO1    => OPEN,
    CO2    => OPEN,
    CO3    => OPEN,
    CO4    => OPEN,
    CO5    => OPEN,
    CO6    => OPEN,
    DSRSTI => '0',
    DDRSTI => '0',
    DSRSTO => OPEN,
    DDRSTO => OPEN,
    DI1    => '0',
    DI2    => '0',
    DI3    => '0',
    DI4    => '0',
    DI5    => '0',
    DI6    => '0',
    DO1    => OPEN,
    DO2    => OPEN,
    DO3    => OPEN,
    DO4    => OPEN,
    DO5    => OPEN,
    DO6    => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U_GRAY2BIN definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CDC_U_GRAY2BIN is
port (
    AI : in  std_logic_vector(5 downto 0);
    AO : out std_logic_vector(5 downto 0);
    BI : in  std_logic_vector(5 downto 0);
    BO : out std_logic_vector(5 downto 0)
);
end NX_CDC_U_GRAY2BIN;

architecture NX_RTL of NX_CDC_U_GRAY2BIN is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 4, -- 4: gray2bin
    ck0_edge       => '0',
    ck1_edge       => '0',
    ack_sel        => '0',
    bck_sel        => '0',
    cck_sel        => '0',
    dck_sel        => '0',
    use_asrc_arst  => '0',
    use_adest_arst => '0',
    use_bsrc_arst  => '0',
    use_bdest_arst => '0',
    use_csrc_arst  => '0',
    use_cdest_arst => '0',
    use_dsrc_arst  => '0',
    use_ddest_arst => '0',
    link_BA        => '0',
    link_CB        => '0',
    link_DC        => '0'
)
port map (
    CK1    => '0',
    CK2    => '0',
    ASRSTI => '0',
    ADRSTI => '0',
    ASRSTO => OPEN,
    ADRSTO => OPEN,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => '0',
    BDRSTI => '0',
    BSRSTO => OPEN,
    BDRSTO => OPEN,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => '0',
    CDRSTI => '0',
    CSRSTO => OPEN,
    CDRSTO => OPEN,
    CI1    => '0',
    CI2    => '0',
    CI3    => '0',
    CI4    => '0',
    CI5    => '0',
    CI6    => '0',
    CO1    => OPEN,
    CO2    => OPEN,
    CO3    => OPEN,
    CO4    => OPEN,
    CO5    => OPEN,
    CO6    => OPEN,
    DSRSTI => '0',
    DDRSTI => '0',
    DSRSTO => OPEN,
    DDRSTO => OPEN,
    DI1    => '0',
    DI2    => '0',
    DI3    => '0',
    DI4    => '0',
    DI5    => '0',
    DI6    => '0',
    DO1    => OPEN,
    DO2    => OPEN,
    DO3    => OPEN,
    DO4    => OPEN,
    DO5    => OPEN,
    DO6    => OPEN
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_XCDC_U definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XCDC_U is
generic (
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI     : in  std_logic_vector(5 downto 0);
    AO     : out std_logic_vector(5 downto 0);
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI     : in  std_logic_vector(5 downto 0);
    BO     : out std_logic_vector(5 downto 0);
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI     : in  std_logic_vector(5 downto 0);
    CO     : out std_logic_vector(5 downto 0);
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI     : in  std_logic_vector(5 downto 0);
    DO     : out std_logic_vector(5 downto 0)
);
end NX_XCDC_U;

architecture NX_RTL of NX_XCDC_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_CDC_U
generic (
    mode           : integer := 0;
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end component NX_CDC_U;

begin

cdc: NX_CDC_U
generic map (
    mode           => 5, -- 5: XCDC
    ck0_edge       => ck0_edge,
    ck1_edge       => ck1_edge,
    ack_sel        => ack_sel,
    bck_sel        => bck_sel,
    cck_sel        => cck_sel,
    dck_sel        => dck_sel,
    use_asrc_arst  => use_asrc_arst,
    use_adest_arst => use_adest_arst,
    use_bsrc_arst  => use_bsrc_arst,
    use_bdest_arst => use_bdest_arst,
    use_csrc_arst  => use_csrc_arst,
    use_cdest_arst => use_cdest_arst,
    use_dsrc_arst  => use_dsrc_arst,
    use_ddest_arst => use_ddest_arst,
    link_BA        => link_BA,
    link_CB        => link_CB,
    link_DC        => link_DC
)
port map (
    CK1    => CK1,
    CK2    => CK2,
    ASRSTI => ASRSTI,
    ADRSTI => ADRSTI,
    ASRSTO => ASRSTO,
    ADRSTO => ADRSTO,
    AI1    => AI(0),
    AI2    => AI(1),
    AI3    => AI(2),
    AI4    => AI(3),
    AI5    => AI(4),
    AI6    => AI(5),
    AO1    => AO(0),
    AO2    => AO(1),
    AO3    => AO(2),
    AO4    => AO(3),
    AO5    => AO(4),
    AO6    => AO(5),
    BSRSTI => BSRSTI,
    BDRSTI => BDRSTI,
    BSRSTO => BSRSTO,
    BDRSTO => BDRSTO,
    BI1    => BI(0),
    BI2    => BI(1),
    BI3    => BI(2),
    BI4    => BI(3),
    BI5    => BI(4),
    BI6    => BI(5),
    BO1    => BO(0),
    BO2    => BO(1),
    BO3    => BO(2),
    BO4    => BO(3),
    BO5    => BO(4),
    BO6    => BO(5),
    CSRSTI => CSRSTI,
    CDRSTI => CDRSTI,
    CSRSTO => CSRSTO,
    CDRSTO => CDRSTO,
    CI1    => CI(0),
    CI2    => CI(1),
    CI3    => CI(2),
    CI4    => CI(3),
    CI5    => CI(4),
    CI6    => CI(5),
    CO1    => CO(0),
    CO2    => CO(1),
    CO3    => CO(2),
    CO4    => CO(3),
    CO5    => CO(4),
    CO6    => CO(5),
    DSRSTI => DSRSTI,
    DDRSTI => DDRSTI,
    DSRSTO => DSRSTO,
    DDRSTO => DDRSTO,
    DI1    => DI(0),
    DI2    => DI(1),
    DI3    => DI(2),
    DI4    => DI(3),
    DI5    => DI(4),
    DI6    => DI(5),
    DO1    => DO(0),
    DO2    => DO(1),
    DO3    => DO(2),
    DO4    => DO(3),
    DO5    => DO(4),
    DO6    => DO(5)
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library NX;
use NX.nxPackage.all;

entity NX_CDC_U is
generic (
    mode           : integer := 0; -- 0: 2DFF     
                                   -- 1: 3DFF     
                                   -- 2: bin2gray + 3DFF + gray2bin
                                   -- 3: bin2gray 
                                   -- 4: gray2bin 
                                   -- 5: XCDC
    ck0_edge       : bit := '0';
    ck1_edge       : bit := '0';
    ack_sel        : bit := '0';
    bck_sel        : bit := '0';
    cck_sel        : bit := '0';
    dck_sel        : bit := '0';
    use_asrc_arst  : bit := '0';
    use_adest_arst : bit := '0';
    use_bsrc_arst  : bit := '0';
    use_bdest_arst : bit := '0';
    use_csrc_arst  : bit := '0';
    use_cdest_arst : bit := '0';
    use_dsrc_arst  : bit := '0';
    use_ddest_arst : bit := '0';
    link_BA        : bit := '0';
    link_CB        : bit := '0';
    link_DC        : bit := '0'
);
port (
    CK1    : in  std_logic;
    CK2    : in  std_logic;
    ASRSTI : in  std_logic;
    ADRSTI : in  std_logic;
    ASRSTO : out std_logic;
    ADRSTO : out std_logic;
    AI1    : in  std_logic;
    AI2    : in  std_logic;
    AI3    : in  std_logic;
    AI4    : in  std_logic;
    AI5    : in  std_logic;
    AI6    : in  std_logic;
    AO1    : out std_logic;
    AO2    : out std_logic;
    AO3    : out std_logic;
    AO4    : out std_logic;
    AO5    : out std_logic;
    AO6    : out std_logic;
    BSRSTI : in  std_logic;
    BDRSTI : in  std_logic;
    BSRSTO : out std_logic;
    BDRSTO : out std_logic;
    BI1    : in  std_logic;
    BI2    : in  std_logic;
    BI3    : in  std_logic;
    BI4    : in  std_logic;
    BI5    : in  std_logic;
    BI6    : in  std_logic;
    BO1    : out std_logic;
    BO2    : out std_logic;
    BO3    : out std_logic;
    BO4    : out std_logic;
    BO5    : out std_logic;
    BO6    : out std_logic;
    CSRSTI : in  std_logic;
    CDRSTI : in  std_logic;
    CSRSTO : out std_logic;
    CDRSTO : out std_logic;
    CI1    : in  std_logic;
    CI2    : in  std_logic;
    CI3    : in  std_logic;
    CI4    : in  std_logic;
    CI5    : in  std_logic;
    CI6    : in  std_logic;
    CO1    : out std_logic;
    CO2    : out std_logic;
    CO3    : out std_logic;
    CO4    : out std_logic;
    CO5    : out std_logic;
    CO6    : out std_logic;
    DSRSTI : in  std_logic;
    DDRSTI : in  std_logic;
    DSRSTO : out std_logic;
    DDRSTO : out std_logic;
    DI1    : in  std_logic;
    DI2    : in  std_logic;
    DI3    : in  std_logic;
    DI4    : in  std_logic;
    DI5    : in  std_logic;
    DI6    : in  std_logic;
    DO1    : out std_logic;
    DO2    : out std_logic;
    DO3    : out std_logic;
    DO4    : out std_logic;
    DO5    : out std_logic;
    DO6    : out std_logic
);
end NX_CDC_U;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_CDC_U mode configuration
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use STD.textio.all;
use ieee.std_logic_textio.all;

package regfile_CDC_U_pkg is 
    
    constant cfg_nc_53downto50                       : std_logic_vector( 2 downto 0):=(others => '0');
    constant cfg_nc_45downto40                       : std_logic_vector( 5 downto 0):=(others => '0');
    constant cfg_test_en_i                           : std_logic_vector( 1 downto 0):=(others => '0');
                                                    
    -- DPREG Link Implementation                    
    constant Conf_2_REG_1RW_1RW_DPREG0_DPREG1        : std_logic_vector( 1 to 7 ):="0000000";
    constant Conf_2_REG_1R_1R_SPREG0_SPREG1          : std_logic_vector( 1 to 7 ):="1100000";
    constant Conf_1_REG_1RW_DEEPER                   : std_logic_vector( 1 to 7 ):="0011111";
    constant Conf_1_REG_1RW_WIDER                    : std_logic_vector( 1 to 7 ):="0001101";
    constant Conf_1_REG_2R_1W                        : std_logic_vector( 1 to 7 ):="0001100";

    function cfg_mode ( mode                         : integer; 
                        ck0_edge                     : std_logic;
                        ck1_edge                     : std_logic;
                        ack_sel                      : std_logic;
                        bck_sel                      : std_logic;
                        cck_sel                      : std_logic;
                        dck_sel                      : std_logic;
                        use_asrc_arst                : std_logic;
                        use_adest_arst               : std_logic;    
                        use_bsrc_arst                : std_logic;  
                        use_bdest_arst               : std_logic;   
                        use_csrc_arst                : std_logic;
                        use_cdest_arst               : std_logic;
                        use_dsrc_arst                : std_logic;
                        use_ddest_arst               : std_logic;
                        link_BA                      : std_logic;
                        link_CB                      : std_logic;
                        link_DC                      : std_logic
                        
        ) return std_logic_vector;


end package regfile_CDC_U_pkg;

package body regfile_CDC_U_pkg is 

    function cfg_mode ( mode                         : integer; 
                        ck0_edge                     : std_logic;
                        ck1_edge                     : std_logic;
                        ack_sel                      : std_logic;
                        bck_sel                      : std_logic;
                        cck_sel                      : std_logic;
                        dck_sel                      : std_logic;
                        use_asrc_arst                : std_logic;
                        use_adest_arst               : std_logic;    
                        use_bsrc_arst                : std_logic;  
                        use_bdest_arst               : std_logic;   
                        use_csrc_arst                : std_logic;
                        use_cdest_arst               : std_logic;
                        use_dsrc_arst                : std_logic;
                        use_ddest_arst               : std_logic;
                        link_BA                      : std_logic;
                        link_CB                      : std_logic;
                        link_DC                      : std_logic
                        
        ) return std_logic_vector is
        -- linked
        variable cfg_reg1_wdata_linked_i           : std_logic;
        variable cfg_reg1_waddr_linked_i           : std_logic;
        variable cfg_reg1_raddr_linked_i           : std_logic;
        variable cfg_reg1_cmd_linked_i             : std_logic;
        variable cfg_reg_linked_i                  : std_logic;
            
        --  cfg_reg0  
        variable cfg_reg0_clkrd_inv_i               : std_logic;
        variable cfg_reg0_clkwr_inv_i               : std_logic;
        variable cfg_reg0_cdc_clk_inv_i             : std_logic;
        variable cfg_reg0_spreg_i                   : std_logic;
        variable cfg_reg0_we_all_mask_i             : std_logic;
        variable cfg_reg0_we_mask_i                 : std_logic;
        variable cfg_reg0_addr_mask_i               : std_logic_vector( 4 downto 0);
        variable cfg_reg0_cdc_dpreg_fifo_i          : std_logic;
        variable cfg_reg0_cdc_w2r_arst_dest_sel_i   : std_logic;
        variable cfg_reg0_cdc_w2r_arst_src_sel_i    : std_logic;
        variable cfg_reg0_cdc_w2r_gray_linked_i     : std_logic;
        variable cfg_reg0_cdc_w2r_use_g2b_i         : std_logic;
        variable cfg_reg0_cdc_w2r_use_b2g_i         : std_logic;
        variable cfg_reg0_cdc_w2r_cdc_clk_i         : std_logic;
        variable cfg_reg0_cdc_w2r_use_reg_dest_i    : std_logic;
        variable cfg_reg0_cdc_w2r_use_reg_src_i     : std_logic;
        variable cfg_reg0_cdc_addr_mask_i           : std_logic_vector( 5 downto 0);
        variable cfg_reg0_cdc_r2w_addrd_inv_i       : std_logic_vector( 5 downto 0);
        variable cfg_reg0_cdc_r2w_arst_dest_sel_i   : std_logic;
        variable cfg_reg0_cdc_r2w_arst_src_sel_i    : std_logic;
        variable cfg_reg0_cdc_r2w_gray_linked_i     : std_logic;
        variable cfg_reg0_cdc_r2w_use_g2b_i         : std_logic;
        variable cfg_reg0_cdc_r2w_use_b2g_i         : std_logic;
        variable cfg_reg0_cdc_r2w_cdc_clk_i         : std_logic;
        variable cfg_reg0_cdc_r2w_use_reg_dest_i    : std_logic;
        variable cfg_reg0_cdc_r2w_use_reg_src_i     : std_logic;

        --  cfg_reg1  
        variable cfg_reg1_clkrd_inv_i               : std_logic;
        variable cfg_reg1_clkwr_inv_i               : std_logic;
        variable cfg_reg1_cdc_clk_inv_i             : std_logic;
        variable cfg_reg1_spreg_i                   : std_logic;
        variable cfg_reg1_we_all_mask_i             : std_logic;
        variable cfg_reg1_we_mask_i                 : std_logic;
        variable cfg_reg1_addr_mask_i               : std_logic_vector( 4 downto 0);
        variable cfg_reg1_cdc_dpreg_fifo_i          : std_logic;
        variable cfg_reg1_cdc_w2r_arst_dest_sel_i   : std_logic;
        variable cfg_reg1_cdc_w2r_arst_src_sel_i    : std_logic;
        variable cfg_reg1_cdc_w2r_gray_linked_i     : std_logic;
        variable cfg_reg1_cdc_w2r_use_g2b_i         : std_logic;
        variable cfg_reg1_cdc_w2r_use_b2g_i         : std_logic;
        variable cfg_reg1_cdc_w2r_cdc_clk_i         : std_logic;
        variable cfg_reg1_cdc_w2r_use_reg_dest_i    : std_logic;
        variable cfg_reg1_cdc_w2r_use_reg_src_i     : std_logic;
        variable cfg_reg1_cdc_addr_mask_i           : std_logic_vector( 5 downto 0);
        variable cfg_reg1_cdc_r2w_addrd_inv_i       : std_logic_vector( 5 downto 0);
        variable cfg_reg1_cdc_r2w_arst_dest_sel_i   : std_logic;
        variable cfg_reg1_cdc_r2w_arst_src_sel_i    : std_logic;
       -- variable cfg_reg1_cdc_r2w_gray_linked_i     : std_logic;
        variable cfg_nc_90                          : std_logic;
        variable cfg_reg1_cdc_r2w_use_g2b_i         : std_logic;
        variable cfg_reg1_cdc_r2w_use_b2g_i         : std_logic;
        variable cfg_reg1_cdc_r2w_cdc_clk_i         : std_logic;
        variable cfg_reg1_cdc_r2w_use_reg_dest_i    : std_logic;
        variable cfg_reg1_cdc_r2w_use_reg_src_i     : std_logic;

        variable DPREG_link_implementation          : std_logic_vector(1 to 7);
        
        variable regfile_config                     : std_logic_vector( 95 downto 0);


        begin
        -- mode :
            -- 0: 2DFF      
            -- 1: 3DFF     
            -- 2: bin2gray + 3DFF + gray2bin
            -- 3: bin2gray 
            -- 4: gray2bin 
            -- 5: XCDC

            cfg_reg1_cdc_r2w_use_reg_src_i      := '1' when mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg1_cdc_r2w_use_reg_dest_i     := '1' when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg1_cdc_r2w_use_b2g_i          := '1' when mode = 2 or mode = 3 or mode = 5 else '0';
            cfg_reg1_cdc_r2w_use_g2b_i          := '1' when mode = 2 or mode = 4 or mode = 5 else '0';
            cfg_nc_90                           := '0';
            
            cfg_reg1_cdc_r2w_addrd_inv_i        := "000000";
            cfg_reg1_cdc_addr_mask_i            := "000000";
            cfg_reg1_cdc_w2r_use_reg_dest_i     := '1' when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg1_cdc_w2r_use_reg_src_i      := '1' when mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg1_cdc_w2r_use_b2g_i          := '1' when mode = 2 or mode = 3 or mode = 5 else '0';
            cfg_reg1_cdc_w2r_use_g2b_i          := '1' when mode = 2 or mode = 4 or mode = 5 else '0';
            cfg_reg1_cdc_w2r_gray_linked_i      :=  link_CB when mode = 5 else '0';
            
            cfg_reg1_cdc_dpreg_fifo_i           := '0';
            cfg_reg1_addr_mask_i                := (others => '0'); --cfg_reg1_addr_mask;-- when mode = 1 else "00000";
            cfg_reg1_we_mask_i                  := '0';
            cfg_reg1_we_all_mask_i              := '0';
            
            -- CDC RESET
            cfg_reg1_cdc_w2r_arst_src_sel_i     :=  use_asrc_arst when mode = 1 or mode = 2 else
                                                    use_bsrc_arst when mode = 5 else 
                                                    '0';
                                                    
            cfg_reg1_cdc_w2r_arst_dest_sel_i    := use_adest_arst when mode = 0 or mode = 1 or mode = 2 else
                                                   use_bdest_arst when mode = 5  else
                                                   '0';
            cfg_reg1_cdc_r2w_arst_src_sel_i     := use_bsrc_arst  when mode = 1 or mode = 2 else
                                                   use_dsrc_arst  when mode = 5   else 
                                                   '0';
                                                   
            cfg_reg1_cdc_r2w_arst_dest_sel_i    := use_bdest_arst when mode = 0 or mode = 1 or mode = 2 else
                                                   use_ddest_arst when mode = 5 else
                                                   '0';
            
            cfg_reg0_cdc_w2r_arst_dest_sel_i    := use_adest_arst when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_w2r_arst_src_sel_i     := use_asrc_arst  when mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_r2w_arst_dest_sel_i    := use_bdest_arst when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_r2w_arst_src_sel_i     := use_bsrc_arst  when mode = 1 or mode = 2 or mode = 5 else '0';
            
            
            --cfg_nc_53downto50                   := '0' when mode = 1 else '0';
            --cfg_test_en_i                       := '0' when mode = 1 else '0';
            --cfg_nc_45downto40                   := '0' when mode = 1 else '0';
            
            -- Clock
            cfg_reg1_cdc_r2w_cdc_clk_i          := '0';
            cfg_reg1_cdc_w2r_cdc_clk_i          := ack_sel when mode = 0 or mode = 1 or mode = 2 else
                                                   bck_sel when mode = 5                         else 
                                                   '0';
            
            -- CLK INV
            cfg_reg1_clkwr_inv_i                := '0';
            cfg_reg1_clkrd_inv_i                := '0';
            cfg_reg0_clkrd_inv_i                := '0';
            cfg_reg0_clkwr_inv_i                := '0';
            cfg_reg0_cdc_clk_inv_i              := ck0_edge when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg1_cdc_clk_inv_i              := ck1_edge when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            
            -- -- 0: 2DFF     
               -- 1: 3DFF     
               -- 2: bin2gray + 3DFF + gray2bin
               -- 3: bin2gray 
               -- 4: gray2bin 
               -- 5: XCDC

            DPREG_link_implementation           := -- Conf_2_REG_1R_1W               when mode =  else
                                                    Conf_2_REG_1RW_1RW_DPREG0_DPREG1 when mode = 0 else
                                                    Conf_2_REG_1R_1R_SPREG0_SPREG1   when mode = 1 else
                                                    Conf_1_REG_1RW_DEEPER            when mode = 2 else
                                                    Conf_1_REG_1RW_WIDER             when mode = 3 else
                                                    Conf_1_REG_2R_1W                 when mode = 4 else
                                                    (others => '0');
            
            -- DPREG link implementation
            cfg_reg0_spreg_i                    := '0';
            cfg_reg1_spreg_i                    := '0';
            cfg_reg_linked_i                    := '0';
            cfg_reg1_cmd_linked_i               := '0';
            cfg_reg1_waddr_linked_i             := '0';
            cfg_reg1_wdata_linked_i             := '0';
            cfg_reg1_raddr_linked_i             := '0';
            
            
            cfg_reg0_we_all_mask_i              := '0'; 
            cfg_reg0_we_mask_i                  := '0'; 
            cfg_reg0_addr_mask_i                := "00000";
            cfg_reg0_cdc_dpreg_fifo_i           := '0';
            
            
            cfg_reg0_cdc_w2r_gray_linked_i      :=  link_BA when mode = 5 else '0';
            cfg_reg0_cdc_w2r_use_g2b_i          := '1' when mode = 2 or mode = 4 or mode = 5 else '0';
            cfg_reg0_cdc_w2r_use_b2g_i          := '1' when mode = 2 or mode = 3 or mode = 5 else '0';
            cfg_reg0_cdc_w2r_cdc_clk_i          := ack_sel when mode = 0 or mode = 1 or mode = 2  or mode = 5 else '0';
            cfg_reg0_cdc_w2r_use_reg_dest_i     := '1' when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_w2r_use_reg_src_i      := '1' when mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_addr_mask_i            := "000000";
            cfg_reg0_cdc_r2w_addrd_inv_i        := "000000";
            
            cfg_reg0_cdc_r2w_gray_linked_i      := link_DC when mode = 5 else '0';
            cfg_reg0_cdc_r2w_use_g2b_i          := '1' when mode = 2 or mode = 4 or mode = 5 else '0';
            cfg_reg0_cdc_r2w_use_b2g_i          := '1' when mode = 2 or mode = 3 or mode = 5 else '0';
            cfg_reg0_cdc_r2w_cdc_clk_i          := bck_sel when mode = 0 or mode = 1 or mode = 2  or mode = 5 else '0';
            cfg_reg0_cdc_r2w_use_reg_dest_i     := '1' when mode = 0 or mode = 1 or mode = 2 or mode = 5 else '0';
            cfg_reg0_cdc_r2w_use_reg_src_i      := '1' when mode = 1 or mode = 2 or mode = 5 else '0';

         
            regfile_config(95)               := cfg_reg1_cdc_r2w_use_reg_src_i     ;  
            regfile_config(94)               := cfg_reg1_cdc_r2w_use_reg_dest_i    ;  
            regfile_config(93)               := cfg_reg1_cdc_r2w_cdc_clk_i         ;  
            regfile_config(92)               := cfg_reg1_cdc_r2w_use_b2g_i         ;  
            regfile_config(91)               := cfg_reg1_cdc_r2w_use_g2b_i         ;  
            regfile_config(90)               := cfg_nc_90                          ;  
            regfile_config(89)               := cfg_reg1_cdc_r2w_arst_src_sel_i    ;  
            regfile_config(88)               := cfg_reg1_cdc_r2w_arst_dest_sel_i   ;  
            regfile_config(87 downto 82)     := cfg_reg1_cdc_r2w_addrd_inv_i       ;  
            regfile_config(81 downto 76)     := cfg_reg1_cdc_addr_mask_i           ;  
            regfile_config(75)               := cfg_reg1_cdc_w2r_use_reg_dest_i    ;  
            regfile_config(74)               := cfg_reg1_cdc_w2r_use_reg_src_i     ;  
            regfile_config(73)               := cfg_reg1_cdc_w2r_cdc_clk_i         ;  
            regfile_config(72)               := cfg_reg1_cdc_w2r_use_b2g_i         ;  
            regfile_config(71)               := cfg_reg1_cdc_w2r_use_g2b_i         ;  
            regfile_config(70)               := cfg_reg1_cdc_w2r_gray_linked_i     ;  
            regfile_config(69)               := cfg_reg1_cdc_w2r_arst_src_sel_i    ;  
            regfile_config(68)               := cfg_reg1_cdc_w2r_arst_dest_sel_i   ;  
            regfile_config(67)               := cfg_reg1_cdc_dpreg_fifo_i          ;  
            regfile_config(66 downto 62)     := cfg_reg1_addr_mask_i               ;  
            regfile_config(61)               := cfg_reg1_we_mask_i                 ;  
            regfile_config(60)               := cfg_reg1_we_all_mask_i             ;  
            regfile_config(59)               := cfg_reg1_spreg_i                   ;  
            regfile_config(58)               := cfg_reg1_cdc_clk_inv_i             ;  
            regfile_config(57)               := cfg_reg1_clkwr_inv_i               ;  
            regfile_config(56)               := cfg_reg1_clkrd_inv_i               ;  
            regfile_config(55 downto 53)     := cfg_nc_53downto50                  ;  
            regfile_config(52)               := cfg_reg1_wdata_linked_i            ;  
            regfile_config(51)               := cfg_reg1_waddr_linked_i            ;  
            regfile_config(50)               := cfg_reg1_raddr_linked_i            ;  
            regfile_config(49)               := cfg_reg1_cmd_linked_i              ;  
            regfile_config(48 downto 47)     := cfg_test_en_i                      ;  
            regfile_config(46)               := cfg_reg_linked_i                   ;  
            regfile_config(45 downto 40)     := cfg_nc_45downto40                  ;  
            regfile_config(39)               := cfg_reg0_clkrd_inv_i               ;  
            regfile_config(38)               := cfg_reg0_clkwr_inv_i               ;  
            regfile_config(37)               := cfg_reg0_cdc_clk_inv_i             ;  
            regfile_config(36)               := cfg_reg0_spreg_i                   ;  
            regfile_config(35)               := cfg_reg0_we_all_mask_i             ;  
            regfile_config(34)               := cfg_reg0_we_mask_i                 ;  
            regfile_config(33 downto 29)     := cfg_reg0_addr_mask_i               ;  
            regfile_config(28)               := cfg_reg0_cdc_dpreg_fifo_i          ;  
            regfile_config(27)               := cfg_reg0_cdc_w2r_arst_dest_sel_i   ;  
            regfile_config(26)               := cfg_reg0_cdc_w2r_arst_src_sel_i    ;  
            regfile_config(25)               := cfg_reg0_cdc_w2r_gray_linked_i     ;  
            regfile_config(24)               := cfg_reg0_cdc_w2r_use_g2b_i         ;  
            regfile_config(23)               := cfg_reg0_cdc_w2r_use_b2g_i         ;  
            regfile_config(22)               := cfg_reg0_cdc_w2r_cdc_clk_i         ;  
            regfile_config(21)               := cfg_reg0_cdc_w2r_use_reg_dest_i    ;  
            regfile_config(20)               := cfg_reg0_cdc_w2r_use_reg_src_i     ;  
            regfile_config(19 downto 14)     := cfg_reg0_cdc_addr_mask_i           ;  
            regfile_config(13 downto  8)     := cfg_reg0_cdc_r2w_addrd_inv_i       ;  
            regfile_config( 7)               := cfg_reg0_cdc_r2w_arst_dest_sel_i   ;  
            regfile_config( 6)               := cfg_reg0_cdc_r2w_arst_src_sel_i    ;  
            regfile_config( 5)               := cfg_reg0_cdc_r2w_gray_linked_i     ;  
            regfile_config( 4)               := cfg_reg0_cdc_r2w_use_g2b_i         ;   
            regfile_config( 3)               := cfg_reg0_cdc_r2w_use_b2g_i         ;   
            regfile_config( 2)               := cfg_reg0_cdc_r2w_cdc_clk_i         ;   
            regfile_config( 1)               := cfg_reg0_cdc_r2w_use_reg_dest_i    ;   
            regfile_config( 0)               := cfg_reg0_cdc_r2w_use_reg_src_i     ;  
            
            return regfile_config(95 downto 0);
        
    end cfg_mode;    
    
end package body regfile_CDC_U_pkg;
-- =================================================================================================
--   NX_RFB_U_WRAP definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_RFB_U_WRAP is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK : in  std_logic;
    I   : in  std_logic_vector(17 downto 0);
    O   : out std_logic_vector(17 downto 0);
    RA  : in  std_logic_vector(4 downto 0);
    WA  : in  std_logic_vector(4 downto 0);
    WE  : in  std_logic;
    WEA : in  std_logic
);
end NX_RFB_U_WRAP;

architecture NX_RTL of NX_RFB_U_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

begin

rfb: NX_RFB_U
generic map (
    mode      => 0, -- 0: DPREG
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I(0),
    I2   => I(1),
    I3   => I(2),
    I4   => I(3),
    I5   => I(4),
    I6   => I(5),
    I7   => I(6),
    I8   => I(7),
    I9   => I(8),
    I10  => I(9),
    I11  => I(10),
    I12  => I(11),
    I13  => I(12),
    I14  => I(13),
    I15  => I(14),
    I16  => I(15),
    I17  => I(16),
    I18  => I(17),
    I19  => '0',
    I20  => '0',
    I21  => '0',
    I22  => '0',
    I23  => '0',
    I24  => '0',
    I25  => '0',
    I26  => '0',
    I27  => '0',
    I28  => '0',
    I29  => '0',
    I30  => '0',
    I31  => '0',
    I32  => '0',
    I33  => '0',
    I34  => '0',
    I35  => '0',
    I36  => '0',
    O1   => O(0),
    O2   => O(1),
    O3   => O(2),
    O4   => O(3),
    O5   => O(4),
    O6   => O(5),
    O7   => O(6),
    O8   => O(7),
    O9   => O(8),
    O10  => O(9),
    O11  => O(10),
    O12  => O(11),
    O13  => O(12),
    O14  => O(13),
    O15  => O(14),
    O16  => O(15),
    O17  => O(16),
    O18  => O(17),
    O19  => OPEN,
    O20  => OPEN,
    O21  => OPEN,
    O22  => OPEN,
    O23  => OPEN,
    O24  => OPEN,
    O25  => OPEN,
    O26  => OPEN,
    O27  => OPEN,
    O28  => OPEN,
    O29  => OPEN,
    O30  => OPEN,
    O31  => OPEN,
    O32  => OPEN,
    O33  => OPEN,
    O34  => OPEN,
    O35  => OPEN,
    O36  => OPEN,
    RA1  => RA(0),
    RA2  => RA(1),
    RA3  => RA(2),
    RA4  => RA(3),
    RA5  => RA(4),
    RA6  => '0',
    RA7  => '0',
    RA8  => '0',
    RA9  => '0',
    RA10 => '0',
    WA1  => WA(0),
    WA2  => WA(1),
    WA3  => WA(2),
    WA4  => WA(3),
    WA5  => WA(4),
    WA6  => '0',
    WE   => WE,
    WEA  => WEA
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_RFBSP_U_WRAP definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_RFBSP_U_WRAP is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK : in  std_logic;
    I   : in  std_logic_vector(17 downto 0);
    O   : out std_logic_vector(17 downto 0);
    WA  : in  std_logic_vector(4 downto 0);
    WE  : in  std_logic;
    WEA : in  std_logic
);
end NX_RFBSP_U_WRAP;

architecture NX_RTL of NX_RFBSP_U_WRAP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

begin

rfb: NX_RFB_U
generic map (
    mode      => 1, -- 1: SPREG
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I(0),
    I2   => I(1),
    I3   => I(2),
    I4   => I(3),
    I5   => I(4),
    I6   => I(5),
    I7   => I(6),
    I8   => I(7),
    I9   => I(8),
    I10  => I(9),
    I11  => I(10),
    I12  => I(11),
    I13  => I(12),
    I14  => I(13),
    I15  => I(14),
    I16  => I(15),
    I17  => I(16),
    I18  => I(17),
    I19  => '0',
    I20  => '0',
    I21  => '0',
    I22  => '0',
    I23  => '0',
    I24  => '0',
    I25  => '0',
    I26  => '0',
    I27  => '0',
    I28  => '0',
    I29  => '0',
    I30  => '0',
    I31  => '0',
    I32  => '0',
    I33  => '0',
    I34  => '0',
    I35  => '0',
    I36  => '0',
    O1   => O(0),
    O2   => O(1),
    O3   => O(2),
    O4   => O(3),
    O5   => O(4),
    O6   => O(5),
    O7   => O(6),
    O8   => O(7),
    O9   => O(8),
    O10  => O(9),
    O11  => O(10),
    O12  => O(11),
    O13  => O(12),
    O14  => O(13),
    O15  => O(14),
    O16  => O(15),
    O17  => O(16),
    O18  => O(17),
    O19  => OPEN,
    O20  => OPEN,
    O21  => OPEN,
    O22  => OPEN,
    O23  => OPEN,
    O24  => OPEN,
    O25  => OPEN,
    O26  => OPEN,
    O27  => OPEN,
    O28  => OPEN,
    O29  => OPEN,
    O30  => OPEN,
    O31  => OPEN,
    O32  => OPEN,
    O33  => OPEN,
    O34  => OPEN,
    O35  => OPEN,
    O36  => OPEN,
    RA1  => '0',
    RA2  => '0',
    RA3  => '0',
    RA4  => '0',
    RA5  => '0',
    RA6  => '0',
    RA7  => '0',
    RA8  => '0',
    RA9  => '0',
    RA10 => '0',
    WA1  => WA(0),
    WA2  => WA(1),
    WA3  => WA(2),
    WA4  => WA(3),
    WA5  => WA(4),
    WA6  => '0',
    WE   => WE,
    WEA  => WEA
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_RFB_U definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_RFB_U is
generic (
    mode     : integer := 0; -- 0: DPREG - 1: SPREG - 2: XRF_64x18 - 3: XRF_32x36 - 4: XRF_2R_1W
    wck_edge : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt : string := "" -- memory initial context
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end NX_RFB_U;

----------------------------------------------------------------------------------------------------


----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RFB_U mode configuration
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use STD.textio.all;
use ieee.std_logic_textio.all;

package regfile_U_pkg is 
    
    constant cfg_nc_53downto50                       : std_logic_vector( 2 downto 0):=(others => '0');
    constant cfg_nc_45downto40                       : std_logic_vector( 5 downto 0):=(others => '0');
    constant cfg_test_en_i                           : std_logic_vector( 1 downto 0):=(others => '0');
                                                    
    -- DPREG Link Implementation                    
    constant Conf_2_REG_1RW_1RW_DPREG0_DPREG1        : std_logic_vector( 1 to 7 ):="0000000";
    constant Conf_2_REG_1R_1R_SPREG0_SPREG1          : std_logic_vector( 1 to 7 ):="1100000";
    constant Conf_1_REG_1RW_DEEPER                   : std_logic_vector( 1 to 7 ):="0011111";
    constant Conf_1_REG_1RW_WIDER                    : std_logic_vector( 1 to 7 ):="0001101";
    constant Conf_1_REG_2R_1W                        : std_logic_vector( 1 to 7 ):="0001100";

    function cfg_mode ( mode                         : integer; 
                        cfg_reg1_cdc_r2w_addrd_inv   : std_logic_vector( 5 downto 0);
                        cfg_reg1_cdc_addr_mask       : std_logic_vector( 5 downto 0);
                        cfg_reg1_addr_mask           : std_logic_vector( 4 downto 0);
                        cfg_reg0_addr_mask           : std_logic_vector( 4 downto 0);
                        cfg_reg0_cdc_addr_mask       : std_logic_vector( 5 downto 0);
                        wck_edge                     : std_logic;                      -- 0: write clock rising edge - 1: write clock falling edge
                        cfg_reg0_cdc_r2w_addrd_inv   : std_logic_vector( 5 downto 0)
                        
        ) return std_logic_vector;


end package regfile_U_pkg;

package body regfile_U_pkg is 

    function cfg_mode ( mode                         : integer; 
                        cfg_reg1_cdc_r2w_addrd_inv   : std_logic_vector( 5 downto 0);
                        cfg_reg1_cdc_addr_mask       : std_logic_vector( 5 downto 0);
                        cfg_reg1_addr_mask           : std_logic_vector( 4 downto 0);
                        cfg_reg0_addr_mask           : std_logic_vector( 4 downto 0);
                        cfg_reg0_cdc_addr_mask       : std_logic_vector( 5 downto 0);
                        wck_edge                     : std_logic;                     -- 0: write clock rising edge - 1: write clock falling edge
                        cfg_reg0_cdc_r2w_addrd_inv   : std_logic_vector( 5 downto 0)
                        
        ) return std_logic_vector is
        -- linked
        variable cfg_reg1_wdata_linked_i           : std_logic;
        variable cfg_reg1_waddr_linked_i           : std_logic;
        variable cfg_reg1_raddr_linked_i           : std_logic;
        variable cfg_reg1_cmd_linked_i             : std_logic;
        variable cfg_reg_linked_i                  : std_logic;
            
        --  cfg_reg0  
        variable cfg_reg0_clkrd_inv_i               : std_logic;
        variable cfg_reg0_clkwr_inv_i               : std_logic;
        variable cfg_reg0_cdc_clk_inv_i             : std_logic;
        variable cfg_reg0_spreg_i                   : std_logic;
        variable cfg_reg0_we_all_mask_i             : std_logic;
        variable cfg_reg0_we_mask_i                 : std_logic;
        variable cfg_reg0_addr_mask_i               : std_logic_vector( 4 downto 0);
        variable cfg_reg0_cdc_dpreg_fifo_i          : std_logic;
        variable cfg_reg0_cdc_w2r_arst_dest_sel_i   : std_logic;
        variable cfg_reg0_cdc_w2r_arst_src_sel_i    : std_logic;
        variable cfg_reg0_cdc_w2r_gray_linked_i     : std_logic;
        variable cfg_reg0_cdc_w2r_use_g2b_i         : std_logic;
        variable cfg_reg0_cdc_w2r_use_b2g_i         : std_logic;
        variable cfg_reg0_cdc_w2r_cdc_clk_i         : std_logic;
        variable cfg_reg0_cdc_w2r_use_reg_dest_i    : std_logic;
        variable cfg_reg0_cdc_w2r_use_reg_src_i     : std_logic;
        variable cfg_reg0_cdc_addr_mask_i           : std_logic_vector( 5 downto 0);
        variable cfg_reg0_cdc_r2w_addrd_inv_i       : std_logic_vector( 5 downto 0);
        variable cfg_reg0_cdc_r2w_arst_dest_sel_i   : std_logic;
        variable cfg_reg0_cdc_r2w_arst_src_sel_i    : std_logic;
        variable cfg_reg0_cdc_r2w_gray_linked_i     : std_logic;
        variable cfg_reg0_cdc_r2w_use_g2b_i         : std_logic;
        variable cfg_reg0_cdc_r2w_use_b2g_i         : std_logic;
        variable cfg_reg0_cdc_r2w_cdc_clk_i         : std_logic;
        variable cfg_reg0_cdc_r2w_use_reg_dest_i    : std_logic;
        variable cfg_reg0_cdc_r2w_use_reg_src_i     : std_logic;

        --  cfg_reg1  
        variable cfg_reg1_clkrd_inv_i               : std_logic;
        variable cfg_reg1_clkwr_inv_i               : std_logic;
        variable cfg_reg1_cdc_clk_inv_i             : std_logic;
        variable cfg_reg1_spreg_i                   : std_logic;
        variable cfg_reg1_we_all_mask_i             : std_logic;
        variable cfg_reg1_we_mask_i                 : std_logic;
        variable cfg_reg1_addr_mask_i               : std_logic_vector( 4 downto 0);
        variable cfg_reg1_cdc_dpreg_fifo_i          : std_logic;
        variable cfg_reg1_cdc_w2r_arst_dest_sel_i   : std_logic;
        variable cfg_reg1_cdc_w2r_arst_src_sel_i    : std_logic;
        constant cfg_reg1_cdc_w2r_gray_linked_i     : std_logic:='0'; --nc
        variable cfg_reg1_cdc_w2r_use_g2b_i         : std_logic;
        variable cfg_reg1_cdc_w2r_use_b2g_i         : std_logic;
        variable cfg_reg1_cdc_w2r_cdc_clk_i         : std_logic;
        variable cfg_reg1_cdc_w2r_use_reg_dest_i    : std_logic;
        variable cfg_reg1_cdc_w2r_use_reg_src_i     : std_logic;
        variable cfg_reg1_cdc_addr_mask_i           : std_logic_vector( 5 downto 0);
        variable cfg_reg1_cdc_r2w_addrd_inv_i       : std_logic_vector( 5 downto 0);
        variable cfg_reg1_cdc_r2w_arst_dest_sel_i   : std_logic;
        variable cfg_reg1_cdc_r2w_arst_src_sel_i    : std_logic;
       -- variable cfg_reg1_cdc_r2w_gray_linked_i     : std_logic;
        variable cfg_nc_90                          : std_logic;
        variable cfg_reg1_cdc_r2w_use_g2b_i         : std_logic;
        variable cfg_reg1_cdc_r2w_use_b2g_i         : std_logic;
        variable cfg_reg1_cdc_r2w_cdc_clk_i         : std_logic;
        variable cfg_reg1_cdc_r2w_use_reg_dest_i    : std_logic;
        variable cfg_reg1_cdc_r2w_use_reg_src_i     : std_logic;

        variable DPREG_link_implementation          : std_logic_vector(1 to 7);
        
        variable regfile_config                     : std_logic_vector( 95 downto 0);


        begin
            --  0  : DPREG0 - 1: SPREG - 2: XRF_64x18 - 3: XRF_32x36 - 4: XRF_2R_1W
            
            cfg_reg1_cdc_r2w_use_reg_src_i      := '0';
            cfg_reg1_cdc_r2w_use_reg_dest_i     := '0';
            cfg_reg1_cdc_r2w_use_b2g_i          := '0';
            cfg_reg1_cdc_r2w_use_g2b_i          := '0';
            cfg_nc_90                           := '0';
            
            cfg_reg1_cdc_r2w_addrd_inv_i        := cfg_reg1_cdc_r2w_addrd_inv_i when mode = 1 else "000000";
            cfg_reg1_cdc_addr_mask_i            := cfg_reg1_cdc_addr_mask       when mode = 1 else "000000";
            cfg_reg1_cdc_w2r_use_reg_dest_i     := '0';
            cfg_reg1_cdc_w2r_use_reg_src_i      := '0';
            cfg_reg1_cdc_w2r_use_b2g_i          := '0';
            cfg_reg1_cdc_w2r_use_g2b_i          := '0';
            --cfg_reg1_cdc_w2r_gray_linked_i      := '0' when mode = 1 else '0';
            
            cfg_reg1_cdc_dpreg_fifo_i           := '0';
            cfg_reg1_addr_mask_i                := cfg_reg1_addr_mask;-- when mode = 1 else "00000";
            cfg_reg1_we_mask_i                  := '0';
            cfg_reg1_we_all_mask_i              := '0';
            
            -- CDC RESET
            cfg_reg1_cdc_w2r_arst_src_sel_i     := '0';
            cfg_reg1_cdc_w2r_arst_dest_sel_i    := '0';
            cfg_reg1_cdc_r2w_arst_src_sel_i     := '0';
            cfg_reg1_cdc_r2w_arst_dest_sel_i    := '0';
            
            cfg_reg0_cdc_w2r_arst_dest_sel_i    := '0';
            cfg_reg0_cdc_w2r_arst_src_sel_i     := '0';
            cfg_reg0_cdc_r2w_arst_dest_sel_i    := '0';
            cfg_reg0_cdc_r2w_arst_src_sel_i     := '0';
            
            
            --cfg_nc_53downto50                   := '0' when mode = 1 else '0';
            --cfg_test_en_i                       := '0' when mode = 1 else '0';
            --cfg_nc_45downto40                   := '0' when mode = 1 else '0';
            
            -- Clock
            cfg_reg1_cdc_r2w_cdc_clk_i          := '0';
            cfg_reg1_cdc_w2r_cdc_clk_i          := '0';
            
            -- CLK INV
            cfg_reg1_clkwr_inv_i                := wck_edge;
            cfg_reg1_clkrd_inv_i                := wck_edge;
            cfg_reg0_clkrd_inv_i                := wck_edge;
            cfg_reg0_clkwr_inv_i                := wck_edge;
            cfg_reg0_cdc_clk_inv_i              := '0';
            cfg_reg1_cdc_clk_inv_i              := '0';
            
            --  0  : DPREG0 - 1: SPREG0 - 2: XRF_64x18 - 3: XRF_32x36 - 4: XRF_2R_1W - 
            DPREG_link_implementation           := -- Conf_2_REG_1R_1W               when mode =  else
                                                    Conf_2_REG_1RW_1RW_DPREG0_DPREG1 when mode = 0 else
                                                    Conf_2_REG_1R_1R_SPREG0_SPREG1   when mode = 1 else
                                                    Conf_1_REG_1RW_DEEPER            when mode = 2 else
                                                    Conf_1_REG_1RW_WIDER             when mode = 3 else
                                                    Conf_1_REG_2R_1W                 when mode = 4 else
                                                    (others => '0');
            
            -- DPREG link implementation
            cfg_reg0_spreg_i                    := DPREG_link_implementation(1);
            cfg_reg1_spreg_i                    := DPREG_link_implementation(2);
            cfg_reg_linked_i                    := DPREG_link_implementation(3);
            cfg_reg1_cmd_linked_i               := DPREG_link_implementation(4);
            cfg_reg1_waddr_linked_i             := DPREG_link_implementation(5);
            cfg_reg1_wdata_linked_i             := DPREG_link_implementation(6);
            cfg_reg1_raddr_linked_i             := DPREG_link_implementation(7);
            
            
            cfg_reg0_we_all_mask_i              := '0'; --'1' when mode = 10  else '0';
            cfg_reg0_we_mask_i                  := '0'; --'1' when mode = 10  else '0';
            cfg_reg0_addr_mask_i                := cfg_reg0_addr_mask when mode = 1 else "00000";
            cfg_reg0_cdc_dpreg_fifo_i           := '0';
            
            
            cfg_reg0_cdc_w2r_gray_linked_i      := '0';
            cfg_reg0_cdc_w2r_use_g2b_i          := '0';
            cfg_reg0_cdc_w2r_use_b2g_i          := '0';
            cfg_reg0_cdc_w2r_cdc_clk_i          := '0';
            cfg_reg0_cdc_w2r_use_reg_dest_i     := '0';
            cfg_reg0_cdc_w2r_use_reg_src_i      := '0';
            cfg_reg0_cdc_addr_mask_i            := cfg_reg0_cdc_addr_mask      when mode = 1 else "000000";
            cfg_reg0_cdc_r2w_addrd_inv_i        := cfg_reg0_cdc_r2w_addrd_inv  when mode = 1 else "000000";
            
            cfg_reg0_cdc_r2w_gray_linked_i      := '0';
            cfg_reg0_cdc_r2w_use_g2b_i          := '0';
            cfg_reg0_cdc_r2w_use_b2g_i          := '0';
            cfg_reg0_cdc_r2w_cdc_clk_i          := '0';
            cfg_reg0_cdc_r2w_use_reg_dest_i     := '0';
            cfg_reg0_cdc_r2w_use_reg_src_i      := '0';

         
        regfile_config(95)               := cfg_reg1_cdc_r2w_use_reg_src_i     ;  
        regfile_config(94)               := cfg_reg1_cdc_r2w_use_reg_dest_i    ;  
        regfile_config(93)               := cfg_reg1_cdc_r2w_cdc_clk_i         ;  
        regfile_config(92)               := cfg_reg1_cdc_r2w_use_b2g_i         ;  
        regfile_config(91)               := cfg_reg1_cdc_r2w_use_g2b_i         ;  
        regfile_config(90)               := cfg_nc_90                          ;  
        regfile_config(89)               := cfg_reg1_cdc_r2w_arst_src_sel_i    ;  
        regfile_config(88)               := cfg_reg1_cdc_r2w_arst_dest_sel_i   ;  
        regfile_config(87 downto 82)     := cfg_reg1_cdc_r2w_addrd_inv_i       ;  
        regfile_config(81 downto 76)     := cfg_reg1_cdc_addr_mask_i           ;  
        regfile_config(75)               := cfg_reg1_cdc_w2r_use_reg_dest_i    ;  
        regfile_config(74)               := cfg_reg1_cdc_w2r_use_reg_src_i     ;  
        regfile_config(73)               := cfg_reg1_cdc_w2r_cdc_clk_i         ;  
        regfile_config(72)               := cfg_reg1_cdc_w2r_use_b2g_i         ;  
        regfile_config(71)               := cfg_reg1_cdc_w2r_use_g2b_i         ;  
        regfile_config(70)               := cfg_reg1_cdc_w2r_gray_linked_i     ;  
        regfile_config(69)               := cfg_reg1_cdc_w2r_arst_src_sel_i    ;  
        regfile_config(68)               := cfg_reg1_cdc_w2r_arst_dest_sel_i   ;  
        regfile_config(67)               := cfg_reg1_cdc_dpreg_fifo_i          ;  
        regfile_config(66 downto 62)     := cfg_reg1_addr_mask_i               ;  
        regfile_config(61)               := cfg_reg1_we_mask_i                 ;  
        regfile_config(60)               := cfg_reg1_we_all_mask_i             ;  
        regfile_config(59)               := cfg_reg1_spreg_i                   ;  
        regfile_config(58)               := cfg_reg1_cdc_clk_inv_i             ;  
        regfile_config(57)               := cfg_reg1_clkwr_inv_i               ;  
        regfile_config(56)               := cfg_reg1_clkrd_inv_i               ;  
        regfile_config(55 downto 53)     := cfg_nc_53downto50                  ;  
        regfile_config(52)               := cfg_reg1_wdata_linked_i            ;  
        regfile_config(51)               := cfg_reg1_waddr_linked_i            ;  
        regfile_config(50)               := cfg_reg1_raddr_linked_i            ;  
        regfile_config(49)               := cfg_reg1_cmd_linked_i              ;  
        regfile_config(48 downto 47)     := cfg_test_en_i                      ;  
        regfile_config(46)               := cfg_reg_linked_i                   ;  
        regfile_config(45 downto 40)     := cfg_nc_45downto40                  ;  
        regfile_config(39)               := cfg_reg0_clkrd_inv_i               ;  
        regfile_config(38)               := cfg_reg0_clkwr_inv_i               ;  
        regfile_config(37)               := cfg_reg0_cdc_clk_inv_i             ;  
        regfile_config(36)               := cfg_reg0_spreg_i                   ;  
        regfile_config(35)               := cfg_reg0_we_all_mask_i             ;  
        regfile_config(34)               := cfg_reg0_we_mask_i                 ;  
        regfile_config(33 downto 29)     := cfg_reg0_addr_mask_i               ;  
        regfile_config(28)               := cfg_reg0_cdc_dpreg_fifo_i          ;  
        regfile_config(27)               := cfg_reg0_cdc_w2r_arst_dest_sel_i   ;  
        regfile_config(26)               := cfg_reg0_cdc_w2r_arst_src_sel_i    ;  
        regfile_config(25)               := cfg_reg0_cdc_w2r_gray_linked_i     ;  
        regfile_config(24)               := cfg_reg0_cdc_w2r_use_g2b_i         ;  
        regfile_config(23)               := cfg_reg0_cdc_w2r_use_b2g_i         ;  
        regfile_config(22)               := cfg_reg0_cdc_w2r_cdc_clk_i         ;  
        regfile_config(21)               := cfg_reg0_cdc_w2r_use_reg_dest_i    ;  
        regfile_config(20)               := cfg_reg0_cdc_w2r_use_reg_src_i     ;  
        regfile_config(19 downto 14)     := cfg_reg0_cdc_addr_mask_i           ;  
        regfile_config(13 downto  8)     := cfg_reg0_cdc_r2w_addrd_inv_i       ;  
        regfile_config( 7)               := cfg_reg0_cdc_r2w_arst_dest_sel_i   ;  
        regfile_config( 6)               := cfg_reg0_cdc_r2w_arst_src_sel_i    ;  
        regfile_config( 5)               := cfg_reg0_cdc_r2w_gray_linked_i     ;  
        regfile_config( 4)               := cfg_reg0_cdc_r2w_use_g2b_i         ;   
        regfile_config( 3)               := cfg_reg0_cdc_r2w_use_b2g_i         ;   
        regfile_config( 2)               := cfg_reg0_cdc_r2w_cdc_clk_i         ;   
        regfile_config( 1)               := cfg_reg0_cdc_r2w_use_reg_dest_i    ;   
        regfile_config( 0)               := cfg_reg0_cdc_r2w_use_reg_src_i     ;  
        
        return regfile_config(95 downto 0);
        
    end cfg_mode;    
    
end package body regfile_U_pkg;
-- =================================================================================================
--   NX_XRFB_64x18 definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XRFB_64x18 is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK : in  std_logic;
    I   : in  std_logic_vector(17 downto 0);
    O   : out std_logic_vector(17 downto 0);
    RA  : in  std_logic_vector(5 downto 0);
    WA  : in  std_logic_vector(5 downto 0);
    WE  : in  std_logic;
    WEA : in  std_logic
);
end NX_XRFB_64x18;

architecture NX_RTL of NX_XRFB_64x18 is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

begin

rfb: NX_RFB_U
generic map (
    mode      => 2, -- 2: DPREG_64x18
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I(0),
    I2   => I(1),
    I3   => I(2),
    I4   => I(3),
    I5   => I(4),
    I6   => I(5),
    I7   => I(6),
    I8   => I(7),
    I9   => I(8),
    I10  => I(9),
    I11  => I(10),
    I12  => I(11),
    I13  => I(12),
    I14  => I(13),
    I15  => I(14),
    I16  => I(15),
    I17  => I(16),
    I18  => I(17),
    I19  => '0',
    I20  => '0',
    I21  => '0',
    I22  => '0',
    I23  => '0',
    I24  => '0',
    I25  => '0',
    I26  => '0',
    I27  => '0',
    I28  => '0',
    I29  => '0',
    I30  => '0',
    I31  => '0',
    I32  => '0',
    I33  => '0',
    I34  => '0',
    I35  => '0',
    I36  => '0',
    O1   => O(0),
    O2   => O(1),
    O3   => O(2),
    O4   => O(3),
    O5   => O(4),
    O6   => O(5),
    O7   => O(6),
    O8   => O(7),
    O9   => O(8),
    O10  => O(9),
    O11  => O(10),
    O12  => O(11),
    O13  => O(12),
    O14  => O(13),
    O15  => O(14),
    O16  => O(15),
    O17  => O(16),
    O18  => O(17),
    O19  => OPEN,
    O20  => OPEN,
    O21  => OPEN,
    O22  => OPEN,
    O23  => OPEN,
    O24  => OPEN,
    O25  => OPEN,
    O26  => OPEN,
    O27  => OPEN,
    O28  => OPEN,
    O29  => OPEN,
    O30  => OPEN,
    O31  => OPEN,
    O32  => OPEN,
    O33  => OPEN,
    O34  => OPEN,
    O35  => OPEN,
    O36  => OPEN,
    RA1  => RA(0),
    RA2  => RA(1),
    RA3  => RA(2),
    RA4  => RA(3),
    RA5  => RA(4),
    RA6  => RA(5),
    RA7  => '0',
    RA8  => '0',
    RA9  => '0',
    RA10 => '0',
    WA1  => WA(0),
    WA2  => WA(1),
    WA3  => WA(2),
    WA4  => WA(3),
    WA5  => WA(4),
    WA6  => WA(5),
    WE   => WE,
    WEA  => WEA
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_XRFB_32x36 definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XRFB_32x36 is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK : in  std_logic;
    I   : in  std_logic_vector(35 downto 0);
    O   : out std_logic_vector(35 downto 0);
    RA  : in  std_logic_vector(4 downto 0);
    WA  : in  std_logic_vector(4 downto 0);
    WE  : in  std_logic;
    WEA : in  std_logic
);
end NX_XRFB_32x36;

architecture NX_RTL of NX_XRFB_32x36 is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

begin

rfb: NX_RFB_U
generic map (
    mode      => 3, -- 3: XRF_32x36
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I(0),
    I2   => I(1),
    I3   => I(2),
    I4   => I(3),
    I5   => I(4),
    I6   => I(5),
    I7   => I(6),
    I8   => I(7),
    I9   => I(8),
    I10  => I(9),
    I11  => I(10),
    I12  => I(11),
    I13  => I(12),
    I14  => I(13),
    I15  => I(14),
    I16  => I(15),
    I17  => I(16),
    I18  => I(17),
    I19  => I(18),
    I20  => I(19),
    I21  => I(20),
    I22  => I(21),
    I23  => I(22),
    I24  => I(23),
    I25  => I(24),
    I26  => I(25),
    I27  => I(26),
    I28  => I(27),
    I29  => I(28),
    I30  => I(29),
    I31  => I(30),
    I32  => I(31),
    I33  => I(32),
    I34  => I(33),
    I35  => I(34),
    I36  => I(35),
    O1   => O(0),
    O2   => O(1),
    O3   => O(2),
    O4   => O(3),
    O5   => O(4),
    O6   => O(5),
    O7   => O(6),
    O8   => O(7),
    O9   => O(8),
    O10  => O(9),
    O11  => O(10),
    O12  => O(11),
    O13  => O(12),
    O14  => O(13),
    O15  => O(14),
    O16  => O(15),
    O17  => O(16),
    O18  => O(17),
    O19  => O(18),
    O20  => O(19),
    O21  => O(20),
    O22  => O(21),
    O23  => O(22),
    O24  => O(23),
    O25  => O(24),
    O26  => O(25),
    O27  => O(26),
    O28  => O(27),
    O29  => O(28),
    O30  => O(29),
    O31  => O(30),
    O32  => O(31),
    O33  => O(32),
    O34  => O(33),
    O35  => O(34),
    O36  => O(35),
    RA1  => RA(0),
    RA2  => RA(1),
    RA3  => RA(2),
    RA4  => RA(3),
    RA5  => RA(4),
    RA6  => '0',
    RA7  => '0',
    RA8  => '0',
    RA9  => '0',
    RA10 => '0',
    WA1 => WA(0),
    WA2 => WA(1),
    WA3 => WA(2),
    WA4 => WA(3),
    WA5 => WA(4),
    WA6 => '0',
    WE  => WE,
    WEA => WEA
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_XRFB_2R_1W definition
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_XRFB_2R_1W is
generic (
    wck_edge  : bit := '0';   -- 0: write clock rising edge - 1: write clock falling edge
    mem_ctxt  : string := "" -- memory initial context
);
port (
    WCK : in  std_logic;
    I   : in  std_logic_vector(17 downto 0);
    AO  : out std_logic_vector(17 downto 0);
    BO  : out std_logic_vector(17 downto 0);
    ARA : in  std_logic_vector(4 downto 0);
    BRA : in  std_logic_vector(4 downto 0);
    WA  : in  std_logic_vector(4 downto 0);
    WE  : in  std_logic;
    WEA : in  std_logic
);
end NX_XRFB_2R_1W;

architecture NX_RTL of NX_XRFB_2R_1W is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RFB_U
generic (
    mode     : integer := 0;
    wck_edge : bit := '0';
    mem_ctxt : string := ""
);
port (
    WCK  : in  std_logic;
    I1   : in  std_logic;
    I2   : in  std_logic;
    I3   : in  std_logic;
    I4   : in  std_logic;
    I5   : in  std_logic;
    I6   : in  std_logic;
    I7   : in  std_logic;
    I8   : in  std_logic;
    I9   : in  std_logic;
    I10  : in  std_logic;
    I11  : in  std_logic;
    I12  : in  std_logic;
    I13  : in  std_logic;
    I14  : in  std_logic;
    I15  : in  std_logic;
    I16  : in  std_logic;
    I17  : in  std_logic;
    I18  : in  std_logic;
    I19  : in  std_logic;
    I20  : in  std_logic;
    I21  : in  std_logic;
    I22  : in  std_logic;
    I23  : in  std_logic;
    I24  : in  std_logic;
    I25  : in  std_logic;
    I26  : in  std_logic;
    I27  : in  std_logic;
    I28  : in  std_logic;
    I29  : in  std_logic;
    I30  : in  std_logic;
    I31  : in  std_logic;
    I32  : in  std_logic;
    I33  : in  std_logic;
    I34  : in  std_logic;
    I35  : in  std_logic;
    I36  : in  std_logic;
    O1   : out std_logic;
    O2   : out std_logic;
    O3   : out std_logic;
    O4   : out std_logic;
    O5   : out std_logic;
    O6   : out std_logic;
    O7   : out std_logic;
    O8   : out std_logic;
    O9   : out std_logic;
    O10  : out std_logic;
    O11  : out std_logic;
    O12  : out std_logic;
    O13  : out std_logic;
    O14  : out std_logic;
    O15  : out std_logic;
    O16  : out std_logic;
    O17  : out std_logic;
    O18  : out std_logic;
    O19  : out std_logic;
    O20  : out std_logic;
    O21  : out std_logic;
    O22  : out std_logic;
    O23  : out std_logic;
    O24  : out std_logic;
    O25  : out std_logic;
    O26  : out std_logic;
    O27  : out std_logic;
    O28  : out std_logic;
    O29  : out std_logic;
    O30  : out std_logic;
    O31  : out std_logic;
    O32  : out std_logic;
    O33  : out std_logic;
    O34  : out std_logic;
    O35  : out std_logic;
    O36  : out std_logic;
    RA1  : in  std_logic;
    RA2  : in  std_logic;
    RA3  : in  std_logic;
    RA4  : in  std_logic;
    RA5  : in  std_logic;
    RA6  : in  std_logic;
    RA7  : in  std_logic;
    RA8  : in  std_logic;
    RA9  : in  std_logic;
    RA10 : in  std_logic;
    WA1  : in  std_logic;
    WA2  : in  std_logic;
    WA3  : in  std_logic;
    WA4  : in  std_logic;
    WA5  : in  std_logic;
    WA6  : in  std_logic;
    WE   : in  std_logic;
    WEA  : in  std_logic
);
end component NX_RFB_U;

begin

rfb: NX_RFB_U
generic map (
    mode      => 4, -- 4: XRF_2R_1W
    wck_edge  => wck_edge,
    mem_ctxt  => mem_ctxt
)
port map (
    WCK  => WCK,
    I1   => I(0),
    I2   => I(1),
    I3   => I(2),
    I4   => I(3),
    I5   => I(4),
    I6   => I(5),
    I7   => I(6),
    I8   => I(7),
    I9   => I(8),
    I10  => I(9),
    I11  => I(10),
    I12  => I(11),
    I13  => I(12),
    I14  => I(13),
    I15  => I(14),
    I16  => I(15),
    I17  => I(16),
    I18  => I(17),
    I19  => '0',
    I20  => '0',
    I21  => '0',
    I22  => '0',
    I23  => '0',
    I24  => '0',
    I25  => '0',
    I26  => '0',
    I27  => '0',
    I28  => '0',
    I29  => '0',
    I30  => '0',
    I31  => '0',
    I32  => '0',
    I33  => '0',
    I34  => '0',
    I35  => '0',
    I36  => '0',
    O1   => AO(0),
    O2   => AO(1),
    O3   => AO(2),
    O4   => AO(3),
    O5   => AO(4),
    O6   => AO(5),
    O7   => AO(6),
    O8   => AO(7),
    O9   => AO(8),
    O10  => AO(9),
    O11  => AO(10),
    O12  => AO(11),
    O13  => AO(12),
    O14  => AO(13),
    O15  => AO(14),
    O16  => AO(15),
    O17  => AO(16),
    O18  => AO(17),
    O19  => BO(0),
    O20  => BO(1),
    O21  => BO(2),
    O22  => BO(3),
    O23  => BO(4),
    O24  => BO(5),
    O25  => BO(6),
    O26  => BO(7),
    O27  => BO(8),
    O28  => BO(9),
    O29  => BO(10),
    O30  => BO(11),
    O31  => BO(12),
    O32  => BO(13),
    O33  => BO(14),
    O34  => BO(15),
    O35  => BO(16),
    O36  => BO(17),
    RA1  => ARA(0),
    RA2  => ARA(1),
    RA3  => ARA(2),
    RA4  => ARA(3),
    RA5  => ARA(4),
    RA6  => BRA(0),
    RA7  => BRA(1),
    RA8  => BRA(2),
    RA9  => BRA(3),
    RA10 => BRA(4),
    WA1 => WA(0),
    WA2 => WA(1),
    WA3 => WA(2),
    WA4 => WA(3),
    WA5 => WA(4),
    WA6 => '0',
    WE  => WE,
    WEA => WEA
);
end NX_RTL;

----------------------------------------------------------------------------------------------------
-- =================================================================================================
--   NX_SER definition                                                                  2018/10/15
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_SER is
generic (
    data_size            : integer range 2 to 10 := 5;	-- Number of serialization factor
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0") or differential ("1")
    slewRate             : string := "";		-- Slow, Medium or Fast
    outputDelayLine      : string := "";		-- "0_to_63_delay_value"
    outputCapacity       : string := "";		-- 0 to 40 (value in pF)
    -- Delay Control
    spath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay

);
port (
    FCK   : in  std_logic;
    SCK   : in  std_logic;
    R     : in  std_logic;
    I     : in  std_logic_vector(data_size - 1 downto 0);
    IO    : out std_logic;
    -- Delay Control
    DCK   : in std_logic;
    DRL   : in std_logic;
    DS    : in std_logic_vector(1 downto 0);
    DRA   : in std_logic_vector(5 downto 0);
    DRI   : in std_logic_vector(5 downto 0);
    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0)
);
end NX_SER;

-- =================================================================================================
--   NX_DES definition                                                                  2018/10/15
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_DES is
generic (
    data_size            : integer range 2 to 10 := 5;	-- -- Pad location Number of deserialization factor
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0") or differential ("1")
    termination          : string := "";		-- Input impedance adaptatio    terminationReference : string := "";
    terminationReference : string := "";		-- "floating" or "VTT"
    turbo                : string := "";		-- Input impedance adaptation
    weakTermination      : string := "";		-- "floating" or "VTT"
    inputDelayLine       : string := "";		-- "0_to_63_delay_value"
    inputSignalSlope     : string := "";		-- Decimal value "0.5" to "20" (value in V/ns)
    -- Delay Control
    dpath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay

);
port (
    FCK   : in  std_logic;
    SCK   : in  std_logic;
    R     : in  std_logic;
    IO    : in  std_logic;
    O     : out std_logic_vector(data_size - 1 downto 0);
    -- Delay Control
    DCK   : in std_logic;
    DRL   : in std_logic;
    DIG   : in std_logic;
    DS    : in std_logic_vector(1 downto 0);
    DRA   : in std_logic_vector(5 downto 0);
    DRI   : in std_logic_vector(5 downto 0);
    FZ    : in std_logic;
    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0);
    FLD   : out std_logic;
    FLG   : out std_logic
);
end NX_DES;

-- =================================================================================================
--   NX_SERDES definition                                                               2018/10/16
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_SERDES is
generic (
    data_size            : integer range 2 to 10 := 5;	-- Serialiser/deserializer factor 
    location             : string := "";		-- Pad location
    standard             : string := "";		-- Pad electrical standard
    drive                : string := "";		-- Pad electrical drive
    differential         : string := "";		-- Single ended ("0" or differential ("1")
    slewRate             : string := "";		-- Slow, Medium or Fast
    termination          : string := "";		-- Input impedance adaptation
    terminationReference : string := "";		-- "floating" or "VTT"
    turbo                : string := "";		-- "true" or "false"
    weakTermination      : string := "";		-- "PullUp" or "None"
    inputDelayLine       : string := "";		-- "O_to_63_delay_value"
    outputDelayLine      : string := "";		-- "O_to_63_delay_value"
    inputSignalSlope     : string := "";		-- Decimal value "0.5" to "20" (value in V/ns)
    outputCapacity       : string := "";		-- "0" to "40" (value in pF)
    cpath_registered     : bit := '0';			-- Use Register in Enable Path ('1')
    -- Delay Control
    spath_dynamic        : bit := '0';			-- 0: off/fixed delay, 1: dynamic delay
    dpath_dynamic        : bit := '0'			-- 0: off/fixed delay, 1: dynamic delay
);
port (
    FCK   : in    std_logic;
    SCK   : in    std_logic;
    RTX   : in    std_logic;
    RRX   : in    std_logic;
    CI    : in    std_logic;
    CCK   : in    std_logic;
    CL    : in    std_logic;
    CR    : in    std_logic;
    I     : in    std_logic_vector(data_size - 1 downto 0);
    IO    : inout std_logic;
    O     : out   std_logic_vector(data_size - 1 downto 0);
    -- Delay Control
    DCK   : in std_logic;
    DRL   : in std_logic;
    DIG   : in std_logic;
    DS    : in std_logic_vector(1 downto 0);
    DRA   : in std_logic_vector(5 downto 0);
    DRI   : in std_logic_vector(5 downto 0);
    FZ    : in std_logic;
    DRO   : out std_logic_vector(5 downto 0);
    DID   : out std_logic_vector(5 downto 0);
    FLD   : out std_logic;
    FLG   : out std_logic
);
end NX_SERDES;

-- NX_SER#{{{#
----------------------------------------------------------------------------------------------------
architecture NX_RTL of NX_SER is

signal I_pad : std_logic;
signal O_pad : std_logic;
signal C_pad : std_logic;
signal sync  : std_logic;
signal I_int : std_logic_vector(9 downto 0);

function BOOL_TO_STR(X : boolean)
  return string is
begin
  if X then
    return "true";
  else
    return "false";
  end if;
end BOOL_TO_STR;

constant spath_delay_on : string := BOOL_TO_STR((outputDelayLine /= "") or (spath_dynamic = '1'));

attribute syn_noprune : boolean;

begin

-- MEDIUM/LARGE#{{{#
SER_M : if NX_SYMBOL /= "NG_U" generate
-- ML ----------------------------------------------------------------------------------------------

signal LINKN : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
signal LINKP : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

begin

I_net: for j in 0 to (data_size - 1) generate
    I_int(j) <= I(j);
end generate;

I_dummy: for j in data_size to 9 generate
    I_int(j) <= '0';
end generate;

single_ser: if (data_size <= 5) generate
attribute syn_noprune of iodx : label is true;
begin

    iobx: NX_IOB_O generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, outputDelayOn        => spath_delay_on
	, outputDelayLine      => outputDelayLine
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		   port map (I => I_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_M generic map (
		   epath_mode      => b"0100"
		 , cpath_mode      => b"0001"
		 , location        => location
		 , symbol          => "SER"
		 )
		 port map (
			   EI1  => I_int(0)
			 , EI2  => I_int(1)
			 , EI3  => I_int(2)
			 , EI4  => I_int(3)
			 , EI5  => I_int(4)
			 , RI   => OPEN
			 , EO   => I_pad
			 , CO   => C_pad
			 , LINK => LINKP
		);
end generate;

large_ser: if (5 < data_size) generate
attribute syn_noprune of iodp : label is true;
attribute syn_noprune of iodn : label is true;
begin

    iobp: NX_IOB_O generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, outputDelayOn        => spath_delay_on
	, outputDelayLine      => outputDelayLine
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		   port map (I => I_pad, C => C_pad, IO => IO);

    iodp: NX_IOM_DRIVER_M generic map (
		   epath_init      => '1'
		 , epath_mode      => b"0100"
		 , cpath_mode      => b"0001"
		 , location        => location
		 , symbol          => "SER"
		 )
		 port map (
			    EI1  => I_int(0)
			  , EI2  => I_int(1)
			  , EI3  => I_int(2)
			  , EI4  => I_int(3)
			  , EI5  => I_int(4)
			  , RI   => OPEN
			  , EO   => I_pad
			  , CO   => C_pad
			  , LINK => LINKP
		);

    iodn: NX_IOM_DRIVER_M generic map (
		   epath_init      => '1'
		 , epath_mode      => b"0100"
		 , cpath_mode      => b"0001"
		 , chained         => '1'
		 , symbol          => "SER_C"
		 )
		 port map (
			    EI1  => I_int(5)
			  , EI2  => I_int(6)
			  , EI3  => I_int(7)
			  , EI4  => I_int(8)
			  , EI5  => I_int(9)
			  , RI   => OPEN
			  , EO   => OPEN
			  , CO   => OPEN
			  , LINK => LINKN
		);
end generate;

iom: NX_IOM_SERDES_M generic map (data_size => data_size, location => location)
		   port map (
			      RTCK  => FCK	    -- ECK
			    , WTCK  => SCK
			    , TRST  => R	    -- ER
			    , DCK   => DCK
			    , DRL   => DRL
			    , DS    => DS
			    , DRA   => DRA
			    , DRI   => DRI
			    , DRO   => DRO
			    , DID   => DID
			    , LINKN => LINKN
			    , LINKP => LINKP
		   );
-- ML ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

-- ULTRA#{{{#
SER_U : if NX_SYMBOL = "NG_U" generate
-- U  ----------------------------------------------------------------------------------------------

signal LINK  : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

-- EMULATION [[[

signal GVON  : std_logic_vector(2 downto 0);
signal GVIN  : std_logic_vector(2 downto 0);
signal GVDN  : std_logic_vector(2 downto 0);
signal GPA   : std_logic_vector(3 downto 0);

-- EMULATION ]]]

begin

I_net: for j in 0 to (data_size - 1) generate
    I_int(j) <= I(j);
end generate;

I_dummy: for j in data_size to 9 generate
    I_int(j) <= '0';
end generate;

single_ser: if (data_size <= 8) generate
attribute syn_noprune of iodx : label is true;
begin

    iobx: NX_IOB_O generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, outputDelayOn        => spath_delay_on
	, outputDelayLine      => outputDelayLine
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		   port map (I => I_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_U generic map (
		   epath_mode      => b"0100"
		 , cpath_mode      => b"0001"
		 , location        => location
		 , symbol          => "SER"
		 )
		 port map (
			   EI1  => I_int(0)
			 , EI2  => I_int(1)
			 , EI3  => I_int(2)
			 , EI4  => I_int(3)
			 , EI5  => I_int(4)
			 , EI6  => I_int(5)
			 , EI7  => I_int(6)
			 , EI8  => I_int(7)
			 , RI   => OPEN
			 , EO   => I_pad
			 , CO   => C_pad
			 , LINK => LINK
		);
end generate;

large_ser: if (8 < data_size) generate
end generate;

cvt: NX_IOM_BIN2GRP
		   port map (
			      LA   => DRA
			    , GS   => DRL
			    , PA   => GPA
			    , GVON => GVON
			    , GVIN => GVIN
			    , GVDN => GVDN
		   );

iom: NX_IOM_SERDES_U generic map (data_size => data_size, location => location)
		   port map (
			      FCK   => FCK
			    , SCK   => SCK
			--  , LDRN
			--  , DRWDS
			--  , DRWEN
			--  , DRE
			    , DRON  => GVON
			    , DRIN  => GVIN
			    , DRDN  => GVDN
			    , DRA   => GPA
			    , DRI   => DRI
			    , FA    => DRA
			--  , FZ
			--  , ALD
			--  , ALT
			    , DRO   => DRO
			    , DID   => DID
			--  , FLD
			--  , FLG
			    , LINK  => LINK
		   );
-- U  ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

end NX_RTL;
-- #}}}#

-- NX_DES#{{{#
----------------------------------------------------------------------------------------------------
architecture NX_RTL of NX_DES is

signal I_pad : std_logic;
signal O_pad : std_logic;
signal C_pad : std_logic;
signal sync  : std_logic;
signal O_int : std_logic_vector(9 downto 0);

function BOOL_TO_STR(X : boolean)
  return string is
begin
  if X then
    return "true";
  else
    return "false";
  end if;
end BOOL_TO_STR;

constant dpath_delay_on : string := BOOL_TO_STR((inputDelayLine /= "") or (dpath_dynamic = '1'));

begin

-- MEDIUM/LARGE#{{{#
DES_M : if NX_SYMBOL /= "NG_U" generate
-- ML ----------------------------------------------------------------------------------------------

signal LINKN : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
signal LINKP : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

begin

O_net: for j in 0 to (data_size - 1) generate
    O(j) <= O_int(j);
end generate;

single_des: if (data_size <= 5) generate

    iobx: NX_IOB_I generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, inputDelayLine       => inputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, locked               => '1'
    )
		   port map (O => O_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_M generic map (
		   rpath_init      => '1'
		 , rpath_mode      => b"0100"
		 , rpath_dynamic   => dpath_dynamic
		 , cpath_mode      => b"0000"
		 , location        => location
		 , symbol          => "DES_D"
		 )
		 port map (
			    RO1  => O_int(4)
			  , RO2  => O_int(3)
			  , RO3  => O_int(2)
			  , RO4  => O_int(1)
			  , RO5  => O_int(0)
			  , RI   => O_pad
			  , EO   => I_pad
			  , CO   => C_pad
			  , LINK => LINKP
		);
end generate;

large_des: if (5 < data_size) generate

    iobp: NX_IOB_I generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, inputDelayLine       => inputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, locked               => '1'
    )
		   port map (O => O_pad, C => C_pad, IO => IO);

    iodp: NX_IOM_DRIVER_M generic map (
		   rpath_init      => '1'
		 , rpath_mode      => b"0100"
		 , rpath_dynamic   => dpath_dynamic
		 , cpath_mode      => b"0000"
		 , location        => location
		 , symbol          => "DES_D"
		 )
		 port map (
			    RO1  => O_int(9)
			  , RO2  => O_int(8)
			  , RO3  => O_int(7)
			  , RO4  => O_int(6)
			  , RO5  => O_int(5)
			  , RI   => O_pad
			  , EO   => I_pad
			  , CO   => C_pad
			  , LINK => LINKP
		);

    iodn: NX_IOM_DRIVER_M generic map (
		  rpath_init       => '1'
		, rpath_mode       => b"0100"
		, cpath_mode       => b"0000"
		, chained          => '1'
		, symbol           => "DES_DC"
		)
		port map (
			   RO1  => O_int(4)
			 , RO2  => O_int(3)
			 , RO3  => O_int(2)
			 , RO4  => O_int(1)
			 , RO5  => O_int(0)
			 , RI   => OPEN
			 , EO   => OPEN
			 , CO   => OPEN
			 , LINK => LINKN
		);
end generate;

iom: NX_IOM_SERDES_M generic map (data_size => data_size, location => location)
		   port map (
			      RRCK  => SCK
			    , WRCK  => FCK	    -- RCK
			    , RRST  => R	    -- RR
			    , DCK   => DCK
			    , DRL   => DRL
			    , DIG   => DIG
			    , DS    => DS
			    , DRA   => DRA
			    , DRI   => DRI
			    , FZ    => FZ
			    , DRO   => DRO
			    , DID   => DID
			    , FLD   => FLD
			    , FLG   => FLG
			    , LINKN => LINKN
			    , LINKP => LINKP
		   );
-- ML ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

-- ULTRA#{{{#
DES_U : if NX_SYMBOL = "NG_U" generate
-- U  ----------------------------------------------------------------------------------------------

signal LINK  : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

-- EMULATION [[[

signal GVON  : std_logic_vector(2 downto 0);
signal GVIN  : std_logic_vector(2 downto 0);
signal GVDN  : std_logic_vector(2 downto 0);
signal GPA   : std_logic_vector(3 downto 0);

-- EMULATION ]]]

begin

O_net: for j in 0 to (data_size - 1) generate
    O(j) <= O_int(j);
end generate;

single_des: if (data_size <= 8) generate

    iobx: NX_IOB_I generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, inputDelayLine       => inputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, locked               => '1'
    )
		   port map (O => O_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_U generic map (
		   rpath_init      => '1'
		 , rpath_mode      => b"0100"
		 , rpath_dynamic   => dpath_dynamic
		 , cpath_mode      => b"0000"
		 , location        => location
		 , symbol          => "DES_D"
		 )
		 port map (
			    RO1  => O_int(7)
			  , RO2  => O_int(6)
			  , RO3  => O_int(5)
			  , RO4  => O_int(4)
			  , RO5  => O_int(3)
			  , RO6  => O_int(2)
			  , RO7  => O_int(1)
			  , RO8  => O_int(0)
			  , RI   => O_pad
			  , EO   => I_pad
			  , CO   => C_pad
			  , LINK => LINK
		);
end generate;

large_des: if (8 < data_size) generate
end generate;

cvt: NX_IOM_BIN2GRP
		   port map (
			      LA   => DRA
			    , GS   => DRL
			    , PA   => GPA
			    , GVON => GVON
			    , GVIN => GVIN
			    , GVDN => GVDN
		   );

iom: NX_IOM_SERDES_U generic map (data_size => data_size, location => location)
		   port map (
			      FCK   => FCK
			    , SCK   => SCK
			--  , LDRN
			--  , DRWDS
			--  , DRWEN
			--  , DRE
			    , DRON  => GVON
			    , DRIN  => GVIN
			    , DRDN  => GVDN
			    , DRA   => GPA
			    , DRI   => DRI
			    , FA    => DRA
			    , FZ    => FZ
			--  , ALD
			--  , ALT
			    , DRO   => DRO
			    , DID   => DID
			    , FLD   => FLD
			    , FLG   => FLG
			    , LINK  => LINK
		   );
-- U  ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

end NX_RTL;
-- #}}}#

-- NX_SERDES#{{{#
----------------------------------------------------------------------------------------------------
architecture NX_RTL of NX_SERDES is

signal I_pad : std_logic;
signal O_pad : std_logic;
signal C_pad : std_logic;
signal sync  : std_logic;
signal I_int : std_logic_vector(9 downto 0);
signal O_int : std_logic_vector(9 downto 0);

function BOOL_TO_STR(X : boolean)
  return string is
begin
  if X then
    return "true";
  else
    return "false";
  end if;
end BOOL_TO_STR;

type switch_mode is array(bit) of bit_vector(3 downto 0);
constant switch : switch_mode := ('0' => b"0010", '1' => b"0011");
constant cpath_mode : bit_vector(3 downto 0) := switch(cpath_registered);

constant spath_delay_on : string := BOOL_TO_STR((outputDelayLine /= "") or (spath_dynamic = '1'));
constant dpath_delay_on : string := BOOL_TO_STR((inputDelayLine  /= "") or (dpath_dynamic = '1'));

begin

-- MEDIUM/LARGE#{{{#
SERDES_M : if NX_SYMBOL /= "NG_U" generate
-- ML ----------------------------------------------------------------------------------------------

signal LINKN : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);
signal LINKP : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

begin

I_net: for j in 0 to (data_size - 1) generate
    I_int(j) <= I(j);
end generate;

I_dummy: for j in (data_size - 1) to 9 generate
    I_int(j) <= '0';
end generate;

O_net: for j in 0 to (data_size - 1) generate
    O(j) <= O_int(j);
end generate;

single_serdes: if (data_size <= 5) generate

    iobx: NX_IOB generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, outputDelayOn        => spath_delay_on
	, inputDelayLine       => inputDelayLine
	, outputDelayLine      => outputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		 port map (I => I_pad, O => O_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_M generic map (
			       epath_init      => '1'
			     , epath_mode      => b"0100"
			     , rpath_init      => '1'
			     , rpath_mode      => b"0100"
			     , rpath_dynamic   => dpath_dynamic
			     , cpath_mode      => cpath_mode
			     , location        => location
			     , symbol          => "SD_DR"
		)
		port map (
			   EI1  => I_int(0)
			 , EI2  => I_int(1)
			 , EI3  => I_int(2)
			 , EI4  => I_int(3)
			 , EI5  => I_int(4)
			 , RO1  => O_int(4)
			 , RO2  => O_int(3)
			 , RO3  => O_int(2)
			 , RO4  => O_int(1)
			 , RO5  => O_int(0)
			 , CI1  => CI
			 , CL   => CL
			 , CR   => CR
			 , RI   => O_pad
			 , EO   => I_pad
			 , CO   => C_pad
			 , LINK => LINKP
		);
end generate;

large_serdes: if (5 < data_size) generate

    iobp: NX_IOB generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, outputDelayOn        => spath_delay_on
	, inputDelayLine       => inputDelayLine
	, outputDelayLine      => outputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		   port map (I => I_pad, O => O_pad, C => C_pad, IO => IO);

    iodp: NX_IOM_DRIVER_M generic map (
			       epath_init      => '1'
			     , epath_mode      => b"0100"
			     , rpath_init      => '1'
			     , rpath_mode      => b"0100"
			     , rpath_dynamic   => dpath_dynamic
			     , cpath_mode      => cpath_mode
			     , location        => location
			     , symbol          => "SD_DR"
		)
		port map (
			   EI1  => I_int(5)
			 , EI2  => I_int(6)
			 , EI3  => I_int(7)
			 , EI4  => I_int(8)
			 , EI5  => I_int(9)
			 , RO1  => O_int(9)
			 , RO2  => O_int(8)
			 , RO3  => O_int(7)
			 , RO4  => O_int(6)
			 , RO5  => O_int(5)
			 , CI1  => CI
			 , CL   => CL
			 , CR   => CR
			 , RI   => O_pad
			 , EO   => I_pad
			 , CO   => C_pad
			 , LINK => LINKP
		);

    iodn: NX_IOM_DRIVER_M generic map (
			       epath_init      => '1'
			     , epath_mode      => b"0100"
			     , rpath_init      => '1'
			     , rpath_mode      => b"0100"
			     , cpath_mode      => cpath_mode
			     , chained         => '1'
			     , symbol          => "SD_DRC"
		)
		port map (
			   EI1  => I_int(0)
			 , EI2  => I_int(1)
			 , EI3  => I_int(2)
			 , EI4  => I_int(3)
			 , EI5  => I_int(4)
			 , RO1  => O_int(4)
			 , RO2  => O_int(3)
			 , RO3  => O_int(2)
			 , RO4  => O_int(1)
			 , RO5  => O_int(0)
			 , CI1  => CI
			 , CL   => CL
			 , CR   => CR
			 , RI   => OPEN
			 , EO   => OPEN
			 , CO   => OPEN
			 , LINK => LINKN
		);
end generate;

iom: NX_IOM_SERDES_M generic map (data_size => data_size, location => location)
		   port map (
			      RTCK  => FCK	    -- ECK
			    , WTCK  => SCK
			    , RRCK  => SCK
			    , WRCK  => FCK	    -- RCK
			    , TRST  => RTX	    -- ER
			    , RRST  => RRX	    -- RR
			    , CTCK  => CCK	    -- CCK
			    , DCK   => DCK
			    , DRL   => DRL
			    , DIG   => DIG
			    , DS    => DS
			    , DRA   => DRA
			    , DRI   => DRI
			    , FZ    => FZ
			    , DRO   => DRO
			    , DID   => DID
			    , FLD   => FLD
			    , FLG   => FLG
			    , LINKN => LINKN
			    , LINKP => LINKP
		   );
-- ML ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

-- ULTRA#{{{#
SERDES_U : if NX_SYMBOL = "NG_U" generate
-- U  ----------------------------------------------------------------------------------------------

signal LINK  : std_logic_vector(IOM_LINK_SIZE - 1 downto 0);

-- EMULATION [[[

signal GVON  : std_logic_vector(2 downto 0);
signal GVIN  : std_logic_vector(2 downto 0);
signal GVDN  : std_logic_vector(2 downto 0);
signal GPA   : std_logic_vector(3 downto 0);

-- EMULATION ]]]

begin

I_net: for j in 0 to (data_size - 1) generate
    I_int(j) <= I(j);
end generate;

I_dummy: for j in (data_size - 1) to 9 generate
    I_int(j) <= '0';
end generate;

O_net: for j in 0 to (data_size - 1) generate
    O(j) <= O_int(j);
end generate;

single_serdes: if (data_size <= 8) generate

    iobx: NX_IOB generic map (
	  location             => location
	, standard             => standard
	, drive                => drive
	, differential         => differential
	, slewRate             => slewRate
	, termination          => termination
	, terminationReference => terminationReference
	, turbo                => turbo
	, weakTermination      => weakTermination
	, inputDelayOn         => dpath_delay_on
	, outputDelayOn        => spath_delay_on
	, inputDelayLine       => inputDelayLine
	, outputDelayLine      => outputDelayLine
	, inputSignalSlope     => inputSignalSlope
	, outputCapacity       => outputCapacity
	, locked               => '1'
    )
		 port map (I => I_pad, O => O_pad, C => C_pad, IO => IO);

    iodx: NX_IOM_DRIVER_U generic map (
			       epath_init      => '1'
			     , epath_mode      => b"0100"
			     , rpath_init      => '1'
			     , rpath_mode      => b"0100"
			     , rpath_dynamic   => dpath_dynamic
			     , cpath_mode      => cpath_mode
			     , location        => location
			     , symbol          => "SD_DR"
		)
		port map (
			   EI1  => I_int(0)
			 , EI2  => I_int(1)
			 , EI3  => I_int(2)
			 , EI4  => I_int(3)
			 , EI5  => I_int(4)
			 , EI6  => I_int(5)
			 , EI7  => I_int(6)
			 , EI8  => I_int(7)
			 , RO1  => O_int(7)
			 , RO2  => O_int(6)
			 , RO3  => O_int(5)
			 , RO4  => O_int(4)
			 , RO5  => O_int(3)
			 , RO6  => O_int(2)
			 , RO7  => O_int(1)
			 , RO8  => O_int(0)
			 , CI1  => CI
			 , CL   => CL
			 , CR   => CR
			 , RI   => O_pad
			 , EO   => I_pad
			 , CO   => C_pad
			 , LINK => LINK
		);
end generate;

large_serdes: if (8 < data_size) generate
end generate;

cvt: NX_IOM_BIN2GRP
		   port map (
			      LA   => DRA
			    , GS   => DRL
			    , PA   => GPA
			    , GVON => GVON
			    , GVIN => GVIN
			    , GVDN => GVDN
		   );

iom: NX_IOM_SERDES_U generic map (data_size => data_size, location => location)
		   port map (
			      FCK   => FCK
			    , SCK   => SCK
			--  , LDRN
			--  , DRWDS
			--  , DRWEN
			--  , DRE
			    , DRON  => GVON
			    , DRIN  => GVIN
			    , DRDN  => GVDN
			    , DRA   => GPA
			    , DRI   => DRI
			    , FA    => DRA
			    , FZ    => FZ
			--  , ALD
			--  , ALT
			    , DRO   => DRO
			    , DID   => DID
			    , FLD   => FLD
			    , FLG   => FLG
			    , LINK  => LINK
		   );
-- U  ----------------------------------------------------------------------------------------------
end generate;
-- #}}}#

end NX_RTL;
-- #}}}#
-- =================================================================================================
--  NX_SERVICE_U definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_SERVICE_U is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    fabric_otp_user_tst_scanenable_i                         : in std_logic;
    fabric_otp_cfg_loader_read_en_i                          : in std_logic;
    fabric_otp_security_force_pdn1_i                         : in std_logic;
    fabric_otp_security_scanenable_i                         : in std_logic;
    fabric_otp_user_din_i1                                   : in std_logic;
    fabric_otp_user_din_i2                                   : in std_logic;
    fabric_otp_user_din_i3                                   : in std_logic;
    fabric_otp_user_din_i4                                   : in std_logic;
    fabric_otp_user_din_i5                                   : in std_logic;
    fabric_otp_user_din_i6                                   : in std_logic;
    fabric_otp_user_din_i7                                   : in std_logic;
    fabric_otp_user_din_i8                                   : in std_logic;
    fabric_otp_user_din_i9                                   : in std_logic;
    fabric_otp_user_din_i10                                  : in std_logic;
    fabric_otp_user_din_i11                                  : in std_logic;
    fabric_otp_user_din_i12                                  : in std_logic;
    fabric_otp_user_din_i13                                  : in std_logic;
    fabric_otp_user_din_i14                                  : in std_logic;
    fabric_otp_user_din_i15                                  : in std_logic;
    fabric_otp_user_din_i16                                  : in std_logic;
    fabric_otp_user_din_i17                                  : in std_logic;
    fabric_otp_user_din_i18                                  : in std_logic;
    fabric_otp_user_din_i19                                  : in std_logic;
    fabric_otp_user_din_i20                                  : in std_logic;
    fabric_otp_user_din_i21                                  : in std_logic;
    fabric_otp_user_din_i22                                  : in std_logic;
    fabric_otp_user_din_i23                                  : in std_logic;
    fabric_otp_user_din_i24                                  : in std_logic;
    fabric_otp_user_din_i25                                  : in std_logic;
    fabric_otp_user_din_i26                                  : in std_logic;
    fabric_otp_user_din_i27                                  : in std_logic;
    fabric_otp_user_din_i28                                  : in std_logic;
    fabric_otp_user_din_i29                                  : in std_logic;
    fabric_otp_user_din_i30                                  : in std_logic;
    fabric_otp_user_din_i31                                  : in std_logic;
    fabric_otp_user_din_i32                                  : in std_logic;
    fabric_otp_user_din_i33                                  : in std_logic;
    fabric_otp_user_din_i34                                  : in std_logic;
    fabric_otp_user_din_i35                                  : in std_logic;
    fabric_otp_user_din_i36                                  : in std_logic;
    fabric_otp_user_din_i37                                  : in std_logic;
    fabric_otp_user_din_i38                                  : in std_logic;
    fabric_otp_user_din_i39                                  : in std_logic;
    fabric_mrepair_fuse_prgwidth_i1                          : in std_logic;
    fabric_mrepair_fuse_prgwidth_i2                          : in std_logic;
    fabric_mrepair_fuse_prgwidth_i3                          : in std_logic;
    fabric_otp_apb_wdata_i1                                  : in std_logic;
    fabric_otp_apb_wdata_i2                                  : in std_logic;
    fabric_otp_apb_wdata_i3                                  : in std_logic;
    fabric_otp_apb_wdata_i4                                  : in std_logic;
    fabric_otp_apb_wdata_i5                                  : in std_logic;
    fabric_otp_apb_wdata_i6                                  : in std_logic;
    fabric_otp_apb_wdata_i7                                  : in std_logic;
    fabric_otp_apb_wdata_i8                                  : in std_logic;
    fabric_otp_apb_wdata_i9                                  : in std_logic;
    fabric_otp_apb_wdata_i10                                 : in std_logic;
    fabric_otp_apb_wdata_i11                                 : in std_logic;
    fabric_otp_apb_wdata_i12                                 : in std_logic;
    fabric_otp_apb_wdata_i13                                 : in std_logic;
    fabric_otp_apb_wdata_i14                                 : in std_logic;
    fabric_otp_apb_wdata_i15                                 : in std_logic;
    fabric_otp_apb_wdata_i16                                 : in std_logic;
    fabric_otp_apb_wdata_i17                                 : in std_logic;
    fabric_otp_apb_wdata_i18                                 : in std_logic;
    fabric_otp_apb_wdata_i19                                 : in std_logic;
    fabric_otp_apb_wdata_i20                                 : in std_logic;
    fabric_otp_apb_wdata_i21                                 : in std_logic;
    fabric_otp_apb_wdata_i22                                 : in std_logic;
    fabric_otp_apb_wdata_i23                                 : in std_logic;
    fabric_otp_apb_wdata_i24                                 : in std_logic;
    fabric_otp_apb_wdata_i25                                 : in std_logic;
    fabric_otp_apb_wdata_i26                                 : in std_logic;
    fabric_otp_apb_wdata_i27                                 : in std_logic;
    fabric_otp_apb_wdata_i28                                 : in std_logic;
    fabric_otp_apb_wdata_i29                                 : in std_logic;
    fabric_otp_apb_wdata_i30                                 : in std_logic;
    fabric_otp_apb_wdata_i31                                 : in std_logic;
    fabric_otp_apb_wdata_i32                                 : in std_logic;
    fabric_otp_cfg_clk_otpm_disable_i                        : in std_logic;
    fabric_otp_user_disturbcheck_i                           : in std_logic;
    fabric_mrepair_fuse_read_i                               : in std_logic;
    fabric_otp_user_rbact2_i                                 : in std_logic;
    fabric_mrepair_fuse_eccbypass_i                          : in std_logic;
    fabric_otp_user_bistmode_i                               : in std_logic;
    fabric_otp_user_add_i1                                   : in std_logic;
    fabric_otp_user_add_i2                                   : in std_logic;
    fabric_otp_user_add_i3                                   : in std_logic;
    fabric_otp_user_add_i4                                   : in std_logic;
    fabric_otp_user_add_i5                                   : in std_logic;
    fabric_otp_user_add_i6                                   : in std_logic;
    fabric_otp_user_add_i7                                   : in std_logic;
    fabric_otp_user_tm_i                                     : in std_logic;
    fabric_otp_rstn_i                                        : in std_logic;
    fabric_mrepair_fuse_disturbchecked_i                     : in std_logic;
    fabric_otp_user_rbact1_i                                 : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i1                        : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i2                        : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i3                        : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i4                        : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i5                        : in std_logic;
    fabric_parusr_type_i1                                    : in std_logic;
    fabric_parusr_type_i2                                    : in std_logic;
    fabric_mrepair_fuse_redbypass_i                          : in std_logic;
    fabric_otp_user_eccbypass_i                              : in std_logic;
    fabric_otp_user_redbypass_i                              : in std_logic;
    fabric_mrepair_mode_i1                                   : in std_logic;
    fabric_mrepair_mode_i2                                   : in std_logic;
    fabric_mrepair_mode_i3                                   : in std_logic;
    fabric_mrepair_mode_i4                                   : in std_logic;
    fabric_parusr_cs_i                                       : in std_logic;
    fabric_sif_reg_en_i1                                     : in std_logic;
    fabric_sif_reg_en_i2                                     : in std_logic;
    fabric_sif_reg_en_i3                                     : in std_logic;
    fabric_sif_reg_en_i4                                     : in std_logic;
    fabric_sif_reg_en_i5                                     : in std_logic;
    fabric_sif_reg_en_i6                                     : in std_logic;
    fabric_sif_reg_en_i7                                     : in std_logic;
    fabric_sif_reg_en_i8                                     : in std_logic;
    fabric_sif_reg_en_i9                                     : in std_logic;
    fabric_sif_reg_en_i10                                    : in std_logic;
    fabric_sif_reg_en_i11                                    : in std_logic;
    fabric_sif_reg_en_i12                                    : in std_logic;
    fabric_sif_reg_en_i13                                    : in std_logic;
    fabric_sif_reg_en_i14                                    : in std_logic;
    fabric_sif_reg_en_i15                                    : in std_logic;
    fabric_sif_reg_en_i16                                    : in std_logic;
    fabric_sif_reg_en_i17                                    : in std_logic;
    fabric_sif_reg_en_i18                                    : in std_logic;
    fabric_sif_reg_en_i19                                    : in std_logic;
    fabric_sif_reg_en_i20                                    : in std_logic;
    fabric_sif_reg_en_i21                                    : in std_logic;
    fabric_sif_reg_en_i22                                    : in std_logic;
    fabric_sif_reg_en_i23                                    : in std_logic;
    fabric_sif_reg_en_i24                                    : in std_logic;
    fabric_sif_reg_en_i25                                    : in std_logic;
    fabric_sif_reg_en_i26                                    : in std_logic;
    fabric_sif_reg_en_i27                                    : in std_logic;
    fabric_sif_reg_en_i28                                    : in std_logic;
    fabric_sif_reg_en_i29                                    : in std_logic;
    fabric_sif_reg_en_i30                                    : in std_logic;
    fabric_sif_reg_en_i31                                    : in std_logic;
    fabric_sif_reg_en_i32                                    : in std_logic;
    fabric_sif_reg_en_i33                                    : in std_logic;
    fabric_sif_reg_en_i34                                    : in std_logic;
    fabric_sif_reg_en_i35                                    : in std_logic;
    fabric_sif_reg_en_i36                                    : in std_logic;
    fabric_sif_reg_en_i37                                    : in std_logic;
    fabric_sif_reg_en_i38                                    : in std_logic;
    fabric_sif_reg_en_i39                                    : in std_logic;
    fabric_sif_reg_en_i40                                    : in std_logic;
    fabric_sif_reg_en_i41                                    : in std_logic;
    fabric_sif_reg_en_i42                                    : in std_logic;
    fabric_sif_reg_en_i43                                    : in std_logic;
    fabric_sif_reg_en_i44                                    : in std_logic;
    fabric_sif_reg_en_i45                                    : in std_logic;
    fabric_sif_reg_en_i46                                    : in std_logic;
    fabric_sif_reg_en_i47                                    : in std_logic;
    fabric_sif_reg_en_i48                                    : in std_logic;
    fabric_sif_reg_en_i49                                    : in std_logic;
    fabric_sif_reg_en_i50                                    : in std_logic;
    fabric_sif_reg_en_i51                                    : in std_logic;
    fabric_sif_reg_en_i52                                    : in std_logic;
    fabric_sif_reg_en_i53                                    : in std_logic;
    fabric_sif_reg_en_i54                                    : in std_logic;
    fabric_sif_reg_en_i55                                    : in std_logic;
    fabric_sif_reg_en_i56                                    : in std_logic;
    fabric_sif_reg_en_i57                                    : in std_logic;
    fabric_sif_reg_en_i58                                    : in std_logic;
    fabric_sif_reg_en_i59                                    : in std_logic;
    fabric_sif_reg_en_i60                                    : in std_logic;
    fabric_sif_reg_en_i61                                    : in std_logic;
    fabric_sif_reg_en_i62                                    : in std_logic;
    fabric_sif_reg_en_i63                                    : in std_logic;
    fabric_sif_reg_en_i64                                    : in std_logic;
    fabric_sif_reg_en_i65                                    : in std_logic;
    fabric_sif_reg_en_i66                                    : in std_logic;
    fabric_sif_reg_en_i67                                    : in std_logic;
    fabric_sif_reg_en_i68                                    : in std_logic;
    fabric_sif_reg_en_i69                                    : in std_logic;
    fabric_sif_reg_en_i70                                    : in std_logic;
    fabric_sif_reg_en_i71                                    : in std_logic;
    fabric_sif_reg_en_i72                                    : in std_logic;
    fabric_sif_reg_en_i73                                    : in std_logic;
    fabric_sif_reg_en_i74                                    : in std_logic;
    fabric_sif_reg_en_i75                                    : in std_logic;
    fabric_sif_reg_en_i76                                    : in std_logic;
    fabric_sif_reg_en_i77                                    : in std_logic;
    fabric_sif_reg_en_i78                                    : in std_logic;
    fabric_sif_reg_en_i79                                    : in std_logic;
    fabric_sif_reg_en_i80                                    : in std_logic;
    fabric_sif_reg_en_i81                                    : in std_logic;
    fabric_sif_reg_en_i82                                    : in std_logic;
    fabric_sif_reg_en_i83                                    : in std_logic;
    fabric_sif_reg_en_i84                                    : in std_logic;
    fabric_sif_reg_en_i85                                    : in std_logic;
    fabric_sif_reg_en_i86                                    : in std_logic;
    fabric_sif_reg_en_i87                                    : in std_logic;
    fabric_sif_reg_en_i88                                    : in std_logic;
    fabric_sif_reg_en_i89                                    : in std_logic;
    fabric_sif_reg_en_i90                                    : in std_logic;
    fabric_sif_reg_en_i91                                    : in std_logic;
    fabric_sif_reg_en_i92                                    : in std_logic;
    fabric_sif_reg_en_i93                                    : in std_logic;
    fabric_sif_reg_en_i94                                    : in std_logic;
    fabric_sif_reg_en_i95                                    : in std_logic;
    fabric_sif_reg_en_i96                                    : in std_logic;
    fabric_sif_reg_en_i97                                    : in std_logic;
    fabric_sif_reg_en_i98                                    : in std_logic;
    fabric_sif_reg_en_i99                                    : in std_logic;
    fabric_sif_reg_en_i100                                   : in std_logic;
    fabric_sif_reg_en_i101                                   : in std_logic;
    fabric_sif_reg_en_i102                                   : in std_logic;
    fabric_sif_reg_en_i103                                   : in std_logic;
    fabric_sif_reg_en_i104                                   : in std_logic;
    fabric_sif_reg_en_i105                                   : in std_logic;
    fabric_sif_reg_en_i106                                   : in std_logic;
    fabric_sif_reg_en_i107                                   : in std_logic;
    fabric_sif_reg_en_i108                                   : in std_logic;
    fabric_sif_reg_en_i109                                   : in std_logic;
    fabric_sif_reg_en_i110                                   : in std_logic;
    fabric_sif_reg_en_i111                                   : in std_logic;
    fabric_sif_reg_en_i112                                   : in std_logic;
    fabric_sif_reg_en_i113                                   : in std_logic;
    fabric_sif_reg_en_i114                                   : in std_logic;
    fabric_sif_reg_en_i115                                   : in std_logic;
    fabric_sif_reg_en_i116                                   : in std_logic;
    fabric_sif_reg_en_i117                                   : in std_logic;
    fabric_sif_reg_en_i118                                   : in std_logic;
    fabric_sif_reg_en_i119                                   : in std_logic;
    fabric_sif_reg_en_i120                                   : in std_logic;
    fabric_mrepair_fuse_rbact2_i                             : in std_logic;
    fabric_data_from_system_i                                : in std_logic;
    fabric_data_from_bist_i1                                 : in std_logic;
    fabric_data_from_bist_i2                                 : in std_logic;
    fabric_data_from_bist_i3                                 : in std_logic;
    fabric_data_from_bist_i4                                 : in std_logic;
    fabric_data_from_bist_i5                                 : in std_logic;
    fabric_data_from_bist_i6                                 : in std_logic;
    fabric_data_from_bist_i7                                 : in std_logic;
    fabric_data_from_bist_i8                                 : in std_logic;
    fabric_data_from_bist_i9                                 : in std_logic;
    fabric_data_from_bist_i10                                : in std_logic;
    fabric_data_from_bist_i11                                : in std_logic;
    fabric_data_from_bist_i12                                : in std_logic;
    fabric_data_from_bist_i13                                : in std_logic;
    fabric_data_from_bist_i14                                : in std_logic;
    fabric_data_from_bist_i15                                : in std_logic;
    fabric_data_from_bist_i16                                : in std_logic;
    fabric_data_from_bist_i17                                : in std_logic;
    fabric_data_from_bist_i18                                : in std_logic;
    fabric_data_from_bist_i19                                : in std_logic;
    fabric_data_from_bist_i20                                : in std_logic;
    fabric_data_from_bist_i21                                : in std_logic;
    fabric_data_from_bist_i22                                : in std_logic;
    fabric_data_from_bist_i23                                : in std_logic;
    fabric_data_from_bist_i24                                : in std_logic;
    fabric_otp_apb_enable_i                                  : in std_logic;
    fabric_mrepair_fuse_tm_i                                 : in std_logic;
    fabric_otp_security_rbact2_i                             : in std_logic;
    fabric_otp_security_rbact1_i                             : in std_logic;
    fabric_shift_en_i1                                       : in std_logic;
    fabric_shift_en_i2                                       : in std_logic;
    fabric_shift_en_i3                                       : in std_logic;
    fabric_shift_en_i4                                       : in std_logic;
    fabric_shift_en_i5                                       : in std_logic;
    fabric_shift_en_i6                                       : in std_logic;
    fabric_shift_en_i7                                       : in std_logic;
    fabric_shift_en_i8                                       : in std_logic;
    fabric_shift_en_i9                                       : in std_logic;
    fabric_shift_en_i10                                      : in std_logic;
    fabric_shift_en_i11                                      : in std_logic;
    fabric_shift_en_i12                                      : in std_logic;
    fabric_shift_en_i13                                      : in std_logic;
    fabric_shift_en_i14                                      : in std_logic;
    fabric_shift_en_i15                                      : in std_logic;
    fabric_shift_en_i16                                      : in std_logic;
    fabric_shift_en_i17                                      : in std_logic;
    fabric_shift_en_i18                                      : in std_logic;
    fabric_shift_en_i19                                      : in std_logic;
    fabric_shift_en_i20                                      : in std_logic;
    fabric_shift_en_i21                                      : in std_logic;
    fabric_shift_en_i22                                      : in std_logic;
    fabric_shift_en_i23                                      : in std_logic;
    fabric_shift_en_i24                                      : in std_logic;
    fabric_otp_cfg_loader_write_en_i                         : in std_logic;
    fabric_user_data_i1                                      : in std_logic;
    fabric_user_data_i2                                      : in std_logic;
    fabric_user_data_i3                                      : in std_logic;
    fabric_user_data_i4                                      : in std_logic;
    fabric_user_data_i5                                      : in std_logic;
    fabric_user_data_i6                                      : in std_logic;
    fabric_user_data_i7                                      : in std_logic;
    fabric_user_data_i8                                      : in std_logic;
    fabric_user_data_i9                                      : in std_logic;
    fabric_user_data_i10                                     : in std_logic;
    fabric_user_data_i11                                     : in std_logic;
    fabric_user_data_i12                                     : in std_logic;
    fabric_user_data_i13                                     : in std_logic;
    fabric_user_data_i14                                     : in std_logic;
    fabric_user_data_i15                                     : in std_logic;
    fabric_user_data_i16                                     : in std_logic;
    fabric_user_data_i17                                     : in std_logic;
    fabric_user_data_i18                                     : in std_logic;
    fabric_user_data_i19                                     : in std_logic;
    fabric_user_data_i20                                     : in std_logic;
    fabric_user_data_i21                                     : in std_logic;
    fabric_user_data_i22                                     : in std_logic;
    fabric_user_data_i23                                     : in std_logic;
    fabric_user_data_i24                                     : in std_logic;
    fabric_user_data_i25                                     : in std_logic;
    fabric_user_data_i26                                     : in std_logic;
    fabric_user_data_i27                                     : in std_logic;
    fabric_user_data_i28                                     : in std_logic;
    fabric_user_data_i29                                     : in std_logic;
    fabric_user_data_i30                                     : in std_logic;
    fabric_user_data_i31                                     : in std_logic;
    fabric_user_data_i32                                     : in std_logic;
    fabric_mrepair_fuse_suppadd_i                            : in std_logic;
    fabric_mrepair_fuse_prog_i                               : in std_logic;
    fabric_otp_user_wordlock_i                               : in std_logic;
    fabric_ahb_direct_data_i1                                : in std_logic;
    fabric_ahb_direct_data_i2                                : in std_logic;
    fabric_ahb_direct_data_i3                                : in std_logic;
    fabric_ahb_direct_data_i4                                : in std_logic;
    fabric_ahb_direct_data_i5                                : in std_logic;
    fabric_ahb_direct_data_i6                                : in std_logic;
    fabric_ahb_direct_data_i7                                : in std_logic;
    fabric_ahb_direct_data_i8                                : in std_logic;
    fabric_ahb_direct_data_i9                                : in std_logic;
    fabric_ahb_direct_data_i10                               : in std_logic;
    fabric_ahb_direct_data_i11                               : in std_logic;
    fabric_ahb_direct_data_i12                               : in std_logic;
    fabric_ahb_direct_data_i13                               : in std_logic;
    fabric_ahb_direct_data_i14                               : in std_logic;
    fabric_ahb_direct_data_i15                               : in std_logic;
    fabric_ahb_direct_data_i16                               : in std_logic;
    fabric_ahb_direct_data_i17                               : in std_logic;
    fabric_ahb_direct_data_i18                               : in std_logic;
    fabric_ahb_direct_data_i19                               : in std_logic;
    fabric_ahb_direct_data_i20                               : in std_logic;
    fabric_ahb_direct_data_i21                               : in std_logic;
    fabric_ahb_direct_data_i22                               : in std_logic;
    fabric_ahb_direct_data_i23                               : in std_logic;
    fabric_ahb_direct_data_i24                               : in std_logic;
    fabric_ahb_direct_data_i25                               : in std_logic;
    fabric_ahb_direct_data_i26                               : in std_logic;
    fabric_ahb_direct_data_i27                               : in std_logic;
    fabric_ahb_direct_data_i28                               : in std_logic;
    fabric_ahb_direct_data_i29                               : in std_logic;
    fabric_ahb_direct_data_i30                               : in std_logic;
    fabric_ahb_direct_data_i31                               : in std_logic;
    fabric_ahb_direct_data_i32                               : in std_logic;
    fabric_otp_user_prog_i                                   : in std_logic;
    fabric_pd_active_i1                                      : in std_logic;
    fabric_pd_active_i2                                      : in std_logic;
    fabric_pd_active_i3                                      : in std_logic;
    fabric_pd_active_i4                                      : in std_logic;
    fabric_pd_active_i5                                      : in std_logic;
    fabric_pd_active_i6                                      : in std_logic;
    fabric_pd_active_i7                                      : in std_logic;
    fabric_pd_active_i8                                      : in std_logic;
    fabric_pd_active_i9                                      : in std_logic;
    fabric_pd_active_i10                                     : in std_logic;
    fabric_pd_active_i11                                     : in std_logic;
    fabric_pd_active_i12                                     : in std_logic;
    fabric_pd_active_i13                                     : in std_logic;
    fabric_pd_active_i14                                     : in std_logic;
    fabric_pd_active_i15                                     : in std_logic;
    fabric_pd_active_i16                                     : in std_logic;
    fabric_pd_active_i17                                     : in std_logic;
    fabric_pd_active_i18                                     : in std_logic;
    fabric_pd_active_i19                                     : in std_logic;
    fabric_pd_active_i20                                     : in std_logic;
    fabric_pd_active_i21                                     : in std_logic;
    fabric_pd_active_i22                                     : in std_logic;
    fabric_pd_active_i23                                     : in std_logic;
    fabric_pd_active_i24                                     : in std_logic;
    fabric_otp_user_suppadd_i                                : in std_logic;
    fabric_mrepair_fuse_pdn_i                                : in std_logic;
    fabric_otp_security_scanin_i1                            : in std_logic;
    fabric_otp_security_scanin_i2                            : in std_logic;
    fabric_otp_security_scanin_i3                            : in std_logic;
    fabric_otp_security_scanin_i4                            : in std_logic;
    fabric_otp_security_scanin_i5                            : in std_logic;
    fabric_end_encoding_i                                    : in std_logic;
    fabric_jtag_tdo_usr2_i                                   : in std_logic;
    fabric_mrepair_fuse_wordlock_i                           : in std_logic;
    fabric_otp_user_prgwidth_i1                              : in std_logic;
    fabric_otp_user_prgwidth_i2                              : in std_logic;
    fabric_otp_user_prgwidth_i3                              : in std_logic;
    fabric_otp_user_read_i                                   : in std_logic;
    fabric_mrepair_fuse_add_i1                               : in std_logic;
    fabric_mrepair_fuse_add_i2                               : in std_logic;
    fabric_mrepair_fuse_add_i3                               : in std_logic;
    fabric_mrepair_fuse_add_i4                               : in std_logic;
    fabric_mrepair_fuse_add_i5                               : in std_logic;
    fabric_mrepair_fuse_add_i6                               : in std_logic;
    fabric_mrepair_fuse_add_i7                               : in std_logic;
    fabric_mrepair_fuse_bistmode_i                           : in std_logic;
    fabric_jtag_tdo_usr1_i                                   : in std_logic;
    fabric_otp_cfg_clk_fab_en_i                              : in std_logic;
    fabric_io_in_i1                                          : in std_logic;
    fabric_io_in_i2                                          : in std_logic;
    fabric_io_in_i3                                          : in std_logic;
    fabric_io_in_i4                                          : in std_logic;
    fabric_io_in_i5                                          : in std_logic;
    fabric_io_in_i6                                          : in std_logic;
    fabric_io_in_i7                                          : in std_logic;
    fabric_io_in_i8                                          : in std_logic;
    fabric_io_in_i9                                          : in std_logic;
    fabric_io_in_i10                                         : in std_logic;
    fabric_io_in_i11                                         : in std_logic;
    fabric_io_in_i12                                         : in std_logic;
    fabric_io_in_i13                                         : in std_logic;
    fabric_io_in_i14                                         : in std_logic;
    fabric_io_in_i15                                         : in std_logic;
    fabric_io_in_i16                                         : in std_logic;
    fabric_io_in_i17                                         : in std_logic;
    fabric_io_in_i18                                         : in std_logic;
    fabric_io_in_i19                                         : in std_logic;
    fabric_io_in_i20                                         : in std_logic;
    fabric_io_in_i21                                         : in std_logic;
    fabric_io_in_i22                                         : in std_logic;
    fabric_io_in_i23                                         : in std_logic;
    fabric_io_in_i24                                         : in std_logic;
    fabric_io_in_i25                                         : in std_logic;
    fabric_sif_load_en_i1                                    : in std_logic;
    fabric_sif_load_en_i2                                    : in std_logic;
    fabric_sif_load_en_i3                                    : in std_logic;
    fabric_sif_load_en_i4                                    : in std_logic;
    fabric_sif_load_en_i5                                    : in std_logic;
    fabric_sif_load_en_i6                                    : in std_logic;
    fabric_sif_load_en_i7                                    : in std_logic;
    fabric_sif_load_en_i8                                    : in std_logic;
    fabric_sif_load_en_i9                                    : in std_logic;
    fabric_sif_load_en_i10                                   : in std_logic;
    fabric_sif_load_en_i11                                   : in std_logic;
    fabric_sif_load_en_i12                                   : in std_logic;
    fabric_sif_load_en_i13                                   : in std_logic;
    fabric_sif_load_en_i14                                   : in std_logic;
    fabric_sif_load_en_i15                                   : in std_logic;
    fabric_sif_load_en_i16                                   : in std_logic;
    fabric_sif_load_en_i17                                   : in std_logic;
    fabric_sif_load_en_i18                                   : in std_logic;
    fabric_sif_load_en_i19                                   : in std_logic;
    fabric_sif_load_en_i20                                   : in std_logic;
    fabric_sif_load_en_i21                                   : in std_logic;
    fabric_sif_load_en_i22                                   : in std_logic;
    fabric_sif_load_en_i23                                   : in std_logic;
    fabric_sif_load_en_i24                                   : in std_logic;
    fabric_mrepair_fuse_din_i1                               : in std_logic;
    fabric_mrepair_fuse_din_i2                               : in std_logic;
    fabric_mrepair_fuse_din_i3                               : in std_logic;
    fabric_mrepair_fuse_din_i4                               : in std_logic;
    fabric_mrepair_fuse_din_i5                               : in std_logic;
    fabric_mrepair_fuse_din_i6                               : in std_logic;
    fabric_mrepair_fuse_din_i7                               : in std_logic;
    fabric_mrepair_fuse_din_i8                               : in std_logic;
    fabric_mrepair_fuse_din_i9                               : in std_logic;
    fabric_mrepair_fuse_din_i10                              : in std_logic;
    fabric_mrepair_fuse_din_i11                              : in std_logic;
    fabric_mrepair_fuse_din_i12                              : in std_logic;
    fabric_mrepair_fuse_din_i13                              : in std_logic;
    fabric_mrepair_fuse_din_i14                              : in std_logic;
    fabric_mrepair_fuse_din_i15                              : in std_logic;
    fabric_mrepair_fuse_din_i16                              : in std_logic;
    fabric_mrepair_fuse_din_i17                              : in std_logic;
    fabric_mrepair_fuse_din_i18                              : in std_logic;
    fabric_mrepair_fuse_din_i19                              : in std_logic;
    fabric_mrepair_fuse_din_i20                              : in std_logic;
    fabric_mrepair_fuse_din_i21                              : in std_logic;
    fabric_mrepair_fuse_din_i22                              : in std_logic;
    fabric_mrepair_fuse_din_i23                              : in std_logic;
    fabric_mrepair_fuse_din_i24                              : in std_logic;
    fabric_mrepair_fuse_din_i25                              : in std_logic;
    fabric_mrepair_fuse_din_i26                              : in std_logic;
    fabric_mrepair_fuse_din_i27                              : in std_logic;
    fabric_mrepair_fuse_din_i28                              : in std_logic;
    fabric_mrepair_fuse_din_i29                              : in std_logic;
    fabric_mrepair_fuse_din_i30                              : in std_logic;
    fabric_mrepair_fuse_din_i31                              : in std_logic;
    fabric_mrepair_fuse_din_i32                              : in std_logic;
    fabric_mrepair_fuse_din_i33                              : in std_logic;
    fabric_mrepair_fuse_din_i34                              : in std_logic;
    fabric_mrepair_fuse_din_i35                              : in std_logic;
    fabric_mrepair_fuse_din_i36                              : in std_logic;
    fabric_mrepair_fuse_din_i37                              : in std_logic;
    fabric_mrepair_fuse_din_i38                              : in std_logic;
    fabric_mrepair_fuse_din_i39                              : in std_logic;
    fabric_otp_apb_addr_i1                                   : in std_logic;
    fabric_otp_apb_addr_i2                                   : in std_logic;
    fabric_otp_apb_addr_i3                                   : in std_logic;
    fabric_otp_apb_addr_i4                                   : in std_logic;
    fabric_otp_apb_addr_i5                                   : in std_logic;
    fabric_otp_apb_addr_i6                                   : in std_logic;
    fabric_otp_apb_addr_i7                                   : in std_logic;
    fabric_otp_apb_addr_i8                                   : in std_logic;
    fabric_otp_apb_addr_i9                                   : in std_logic;
    fabric_otp_apb_addr_i10                                  : in std_logic;
    fabric_otp_apb_addr_i11                                  : in std_logic;
    fabric_otp_apb_addr_i12                                  : in std_logic;
    fabric_otp_apb_addr_i13                                  : in std_logic;
    fabric_otp_apb_addr_i14                                  : in std_logic;
    fabric_otp_apb_addr_i15                                  : in std_logic;
    fabric_otp_apb_addr_i16                                  : in std_logic;
    fabric_otp_apb_addr_i17                                  : in std_logic;
    fabric_otp_apb_addr_i18                                  : in std_logic;
    fabric_otp_apb_addr_i19                                  : in std_logic;
    fabric_otp_apb_addr_i20                                  : in std_logic;
    fabric_otp_apb_addr_i21                                  : in std_logic;
    fabric_otp_apb_addr_i22                                  : in std_logic;
    fabric_otp_apb_addr_i23                                  : in std_logic;
    fabric_otp_apb_addr_i24                                  : in std_logic;
    fabric_otp_apb_addr_i25                                  : in std_logic;
    fabric_otp_apb_addr_i26                                  : in std_logic;
    fabric_otp_apb_addr_i27                                  : in std_logic;
    fabric_otp_apb_addr_i28                                  : in std_logic;
    fabric_otp_apb_addr_i29                                  : in std_logic;
    fabric_otp_apb_addr_i30                                  : in std_logic;
    fabric_otp_apb_addr_i31                                  : in std_logic;
    fabric_otp_apb_addr_i32                                  : in std_logic;
    fabric_otp_apb_sel_i                                     : in std_logic;
    fabric_mrepair_fuse_rbact1_i                             : in std_logic;
    fabric_mrepair_fuse_configreg_i1                         : in std_logic;
    fabric_mrepair_fuse_configreg_i2                         : in std_logic;
    fabric_mrepair_fuse_configreg_i3                         : in std_logic;
    fabric_mrepair_fuse_configreg_i4                         : in std_logic;
    fabric_mrepair_fuse_configreg_i5                         : in std_logic;
    fabric_mrepair_fuse_configreg_i6                         : in std_logic;
    fabric_mrepair_fuse_configreg_i7                         : in std_logic;
    fabric_mrepair_fuse_configreg_i8                         : in std_logic;
    fabric_mrepair_fuse_configreg_i9                         : in std_logic;
    fabric_mrepair_fuse_configreg_i10                        : in std_logic;
    fabric_mrepair_fuse_configreg_i11                        : in std_logic;
    fabric_mrepair_fuse_configreg_i12                        : in std_logic;
    fabric_mrepair_fuse_configreg_i13                        : in std_logic;
    fabric_mrepair_fuse_configreg_i14                        : in std_logic;
    fabric_mrepair_fuse_configreg_i15                        : in std_logic;
    fabric_mrepair_fuse_configreg_i16                        : in std_logic;
    fabric_mrepair_fuse_configreg_i17                        : in std_logic;
    fabric_mrepair_fuse_configreg_i18                        : in std_logic;
    fabric_mrepair_fuse_configreg_i19                        : in std_logic;
    fabric_mrepair_fuse_configreg_i20                        : in std_logic;
    fabric_mrepair_fuse_configreg_i21                        : in std_logic;
    fabric_mrepair_fuse_configreg_i22                        : in std_logic;
    fabric_mrepair_fuse_configreg_i23                        : in std_logic;
    fabric_mrepair_fuse_configreg_i24                        : in std_logic;
    fabric_mrepair_fuse_configreg_i25                        : in std_logic;
    fabric_mrepair_fuse_configreg_i26                        : in std_logic;
    fabric_mrepair_fuse_configreg_i27                        : in std_logic;
    fabric_mrepair_fuse_configreg_i28                        : in std_logic;
    fabric_mrepair_fuse_configreg_i29                        : in std_logic;
    fabric_mrepair_fuse_configreg_i30                        : in std_logic;
    fabric_mrepair_fuse_configreg_i31                        : in std_logic;
    fabric_mrepair_fuse_configreg_i32                        : in std_logic;
    fabric_otp_cfg_fabric_apb_en_i                           : in std_logic;
    fabric_data_shift_en_i                                   : in std_logic;
    fabric_lowskew_i21                                       : in std_logic;
    fabric_direct_data_i1                                    : in std_logic;
    fabric_direct_data_i2                                    : in std_logic;
    fabric_direct_data_i3                                    : in std_logic;
    fabric_direct_data_i4                                    : in std_logic;
    fabric_direct_data_i5                                    : in std_logic;
    fabric_direct_data_i6                                    : in std_logic;
    fabric_direct_data_i7                                    : in std_logic;
    fabric_direct_data_i8                                    : in std_logic;
    fabric_direct_data_i9                                    : in std_logic;
    fabric_direct_data_i10                                   : in std_logic;
    fabric_direct_data_i11                                   : in std_logic;
    fabric_direct_data_i12                                   : in std_logic;
    fabric_direct_data_i13                                   : in std_logic;
    fabric_direct_data_i14                                   : in std_logic;
    fabric_direct_data_i15                                   : in std_logic;
    fabric_direct_data_i16                                   : in std_logic;
    fabric_direct_data_i17                                   : in std_logic;
    fabric_direct_data_i18                                   : in std_logic;
    fabric_direct_data_i19                                   : in std_logic;
    fabric_direct_data_i20                                   : in std_logic;
    fabric_direct_data_i21                                   : in std_logic;
    fabric_direct_data_i22                                   : in std_logic;
    fabric_direct_data_i23                                   : in std_logic;
    fabric_direct_data_i24                                   : in std_logic;
    fabric_direct_data_i25                                   : in std_logic;
    fabric_direct_data_i26                                   : in std_logic;
    fabric_direct_data_i27                                   : in std_logic;
    fabric_direct_data_i28                                   : in std_logic;
    fabric_direct_data_i29                                   : in std_logic;
    fabric_direct_data_i30                                   : in std_logic;
    fabric_direct_data_i31                                   : in std_logic;
    fabric_direct_data_i32                                   : in std_logic;
    fabric_otp_user_pdn_i                                    : in std_logic;
    fabric_io_oe_i1                                          : in std_logic;
    fabric_io_oe_i2                                          : in std_logic;
    fabric_io_oe_i3                                          : in std_logic;
    fabric_io_oe_i4                                          : in std_logic;
    fabric_io_oe_i5                                          : in std_logic;
    fabric_io_oe_i6                                          : in std_logic;
    fabric_io_oe_i7                                          : in std_logic;
    fabric_io_oe_i8                                          : in std_logic;
    fabric_io_oe_i9                                          : in std_logic;
    fabric_io_oe_i10                                         : in std_logic;
    fabric_io_oe_i11                                         : in std_logic;
    fabric_io_oe_i12                                         : in std_logic;
    fabric_io_oe_i13                                         : in std_logic;
    fabric_io_oe_i14                                         : in std_logic;
    fabric_io_oe_i15                                         : in std_logic;
    fabric_io_oe_i16                                         : in std_logic;
    fabric_io_oe_i17                                         : in std_logic;
    fabric_io_oe_i18                                         : in std_logic;
    fabric_io_oe_i19                                         : in std_logic;
    fabric_io_oe_i20                                         : in std_logic;
    fabric_io_oe_i21                                         : in std_logic;
    fabric_io_oe_i22                                         : in std_logic;
    fabric_io_oe_i23                                         : in std_logic;
    fabric_io_oe_i24                                         : in std_logic;
    fabric_io_oe_i25                                         : in std_logic;
    fabric_parusr_data_i1                                    : in std_logic;
    fabric_parusr_data_i2                                    : in std_logic;
    fabric_parusr_data_i3                                    : in std_logic;
    fabric_parusr_data_i4                                    : in std_logic;
    fabric_parusr_data_i5                                    : in std_logic;
    fabric_parusr_data_i6                                    : in std_logic;
    fabric_parusr_data_i7                                    : in std_logic;
    fabric_parusr_data_i8                                    : in std_logic;
    fabric_parusr_data_i9                                    : in std_logic;
    fabric_parusr_data_i10                                   : in std_logic;
    fabric_parusr_data_i11                                   : in std_logic;
    fabric_parusr_data_i12                                   : in std_logic;
    fabric_parusr_data_i13                                   : in std_logic;
    fabric_parusr_data_i14                                   : in std_logic;
    fabric_parusr_data_i15                                   : in std_logic;
    fabric_parusr_data_i16                                   : in std_logic;
    fabric_otp_apb_write_i                                   : in std_logic;
    fabric_otp_security_testmode_i                           : in std_logic;
    fabric_system_data_to_mem_bist_i1                        : in std_logic;
    fabric_system_data_to_mem_bist_i2                        : in std_logic;
    fabric_system_data_to_mem_bist_i3                        : in std_logic;
    fabric_system_data_to_mem_bist_i4                        : in std_logic;
    fabric_system_data_to_mem_bist_i5                        : in std_logic;
    fabric_system_data_to_mem_bist_i6                        : in std_logic;
    fabric_system_data_to_mem_bist_i7                        : in std_logic;
    fabric_system_data_to_mem_bist_i8                        : in std_logic;
    fabric_system_data_to_mem_bist_i9                        : in std_logic;
    fabric_system_data_to_mem_bist_i10                       : in std_logic;
    fabric_system_data_to_mem_bist_i11                       : in std_logic;
    fabric_system_data_to_mem_bist_i12                       : in std_logic;
    fabric_system_data_to_mem_bist_i13                       : in std_logic;
    fabric_system_data_to_mem_bist_i14                       : in std_logic;
    fabric_system_data_to_mem_bist_i15                       : in std_logic;
    fabric_system_data_to_mem_bist_i16                       : in std_logic;
    fabric_system_data_to_mem_bist_i17                       : in std_logic;
    fabric_system_data_to_mem_bist_i18                       : in std_logic;
    fabric_system_data_to_mem_bist_i19                       : in std_logic;
    fabric_system_data_to_mem_bist_i20                       : in std_logic;
    fabric_system_data_to_mem_bist_i21                       : in std_logic;
    fabric_system_data_to_mem_bist_i22                       : in std_logic;
    fabric_system_data_to_mem_bist_i23                       : in std_logic;
    fabric_system_data_to_mem_bist_i24                       : in std_logic;
    fabric_tst_atpg_mrepair_i                                : in std_logic;
    fabric_mrepair_fuse_tstscanenable_i                      : in std_logic;
    fabric_otp_security_bistmode_i                           : in std_logic;
    fabric_lowskew_i22                                       : in std_logic;
    fabric_lowskew_i23                                       : in std_logic;
    fabric_lowskew_i20                                       : in std_logic;
    fabric_otp_user_configreg_i1                             : in std_logic;
    fabric_otp_user_configreg_i2                             : in std_logic;
    fabric_otp_user_configreg_i3                             : in std_logic;
    fabric_otp_user_configreg_i4                             : in std_logic;
    fabric_otp_user_configreg_i5                             : in std_logic;
    fabric_otp_user_configreg_i6                             : in std_logic;
    fabric_otp_user_configreg_i7                             : in std_logic;
    fabric_otp_user_configreg_i8                             : in std_logic;
    fabric_otp_user_configreg_i9                             : in std_logic;
    fabric_otp_user_configreg_i10                            : in std_logic;
    fabric_otp_user_configreg_i11                            : in std_logic;
    fabric_otp_user_configreg_i12                            : in std_logic;
    fabric_otp_user_configreg_i13                            : in std_logic;
    fabric_otp_user_configreg_i14                            : in std_logic;
    fabric_otp_user_configreg_i15                            : in std_logic;
    fabric_otp_user_configreg_i16                            : in std_logic;
    fabric_otp_user_configreg_i17                            : in std_logic;
    fabric_otp_user_configreg_i18                            : in std_logic;
    fabric_otp_user_configreg_i19                            : in std_logic;
    fabric_otp_user_configreg_i20                            : in std_logic;
    fabric_otp_user_configreg_i21                            : in std_logic;
    fabric_otp_user_configreg_i22                            : in std_logic;
    fabric_otp_user_configreg_i23                            : in std_logic;
    fabric_otp_user_configreg_i24                            : in std_logic;
    fabric_otp_user_configreg_i25                            : in std_logic;
    fabric_otp_user_configreg_i26                            : in std_logic;
    fabric_otp_user_configreg_i27                            : in std_logic;
    fabric_otp_user_configreg_i28                            : in std_logic;
    fabric_otp_user_configreg_i29                            : in std_logic;
    fabric_otp_user_configreg_i30                            : in std_logic;
    fabric_otp_user_configreg_i31                            : in std_logic;
    fabric_otp_user_configreg_i32                            : in std_logic;
    fabric_otp_user_tst_scanin_i1                            : in std_logic;
    fabric_otp_user_tst_scanin_i2                            : in std_logic;
    fabric_otp_user_tst_scanin_i3                            : in std_logic;
    fabric_otp_user_tst_scanin_i4                            : in std_logic;
    fabric_otp_user_tst_scanin_i5                            : in std_logic;
    fabric_sif_update_en_i1                                  : in std_logic;
    fabric_sif_update_en_i2                                  : in std_logic;
    fabric_sif_update_en_i3                                  : in std_logic;
    fabric_sif_update_en_i4                                  : in std_logic;
    fabric_sif_update_en_i5                                  : in std_logic;
    fabric_sif_update_en_i6                                  : in std_logic;
    fabric_sif_update_en_i7                                  : in std_logic;
    fabric_sif_update_en_i8                                  : in std_logic;
    fabric_sif_update_en_i9                                  : in std_logic;
    fabric_sif_update_en_i10                                 : in std_logic;
    fabric_sif_update_en_i11                                 : in std_logic;
    fabric_sif_update_en_i12                                 : in std_logic;
    fabric_sif_update_en_i13                                 : in std_logic;
    fabric_sif_update_en_i14                                 : in std_logic;
    fabric_sif_update_en_i15                                 : in std_logic;
    fabric_sif_update_en_i16                                 : in std_logic;
    fabric_sif_update_en_i17                                 : in std_logic;
    fabric_sif_update_en_i18                                 : in std_logic;
    fabric_sif_update_en_i19                                 : in std_logic;
    fabric_sif_update_en_i20                                 : in std_logic;
    fabric_sif_update_en_i21                                 : in std_logic;
    fabric_sif_update_en_i22                                 : in std_logic;
    fabric_sif_update_en_i23                                 : in std_logic;
    fabric_sif_update_en_i24                                 : in std_logic;
    fabric_mrepair_por_i                                     : in std_logic;
    fabric_mrepair_rst_n_i                                   : in std_logic;
    fabric_mrepair_initn_i                                   : in std_logic;
    fabric_spare_i1                                          : in std_logic;
    fabric_spare_i2                                          : in std_logic;
    fabric_spare_i3                                          : in std_logic;

    fabric_mrepair_fuse_bbad_o                               : out std_logic;
    fabric_jtag_trst_n_o                                     : out std_logic;
    fabric_debug_direct_permission_write_o1                  : out std_logic;
    fabric_debug_direct_permission_write_o2                  : out std_logic;
    fabric_debug_direct_permission_write_o3                  : out std_logic;
    fabric_debug_direct_permission_write_o4                  : out std_logic;
    fabric_otp_security_bist_end1_o                          : out std_logic;
    fabric_parusr_data_val_o                                 : out std_logic;
    fabric_debug_lock_reg_o                                  : out std_logic;
    fabric_debug_security_error_read_o                       : out std_logic;
    fabric_mrepair_fuse_tstscanout_o1                        : out std_logic;
    fabric_mrepair_fuse_tstscanout_o2                        : out std_logic;
    fabric_mrepair_fuse_tstscanout_o3                        : out std_logic;
    fabric_mrepair_fuse_tstscanout_o4                        : out std_logic;
    fabric_mrepair_fuse_tstscanout_o5                        : out std_logic;
    fabric_otp_user_tst_scanout_o1                           : out std_logic;
    fabric_otp_user_tst_scanout_o2                           : out std_logic;
    fabric_otp_user_tst_scanout_o3                           : out std_logic;
    fabric_otp_user_tst_scanout_o4                           : out std_logic;
    fabric_otp_user_tst_scanout_o5                           : out std_logic;
    fabric_sif_update_en_to_bist_o1                          : out std_logic;
    fabric_sif_update_en_to_bist_o2                          : out std_logic;
    fabric_sif_update_en_to_bist_o3                          : out std_logic;
    fabric_sif_update_en_to_bist_o4                          : out std_logic;
    fabric_sif_update_en_to_bist_o5                          : out std_logic;
    fabric_sif_update_en_to_bist_o6                          : out std_logic;
    fabric_sif_update_en_to_bist_o7                          : out std_logic;
    fabric_sif_update_en_to_bist_o8                          : out std_logic;
    fabric_sif_update_en_to_bist_o9                          : out std_logic;
    fabric_sif_update_en_to_bist_o10                         : out std_logic;
    fabric_sif_update_en_to_bist_o11                         : out std_logic;
    fabric_sif_update_en_to_bist_o12                         : out std_logic;
    fabric_sif_update_en_to_bist_o13                         : out std_logic;
    fabric_sif_update_en_to_bist_o14                         : out std_logic;
    fabric_sif_update_en_to_bist_o15                         : out std_logic;
    fabric_sif_update_en_to_bist_o16                         : out std_logic;
    fabric_sif_update_en_to_bist_o17                         : out std_logic;
    fabric_sif_update_en_to_bist_o18                         : out std_logic;
    fabric_sif_update_en_to_bist_o19                         : out std_logic;
    fabric_sif_update_en_to_bist_o20                         : out std_logic;
    fabric_sif_update_en_to_bist_o21                         : out std_logic;
    fabric_sif_update_en_to_bist_o22                         : out std_logic;
    fabric_sif_update_en_to_bist_o23                         : out std_logic;
    fabric_sif_update_en_to_bist_o24                         : out std_logic;
    fabric_otp_user_locked_o                                 : out std_logic;
    fabric_otp_security_bist_bad_o                           : out std_logic;
    fabric_debug_frame_permission_frame_o1                   : out std_logic;
    fabric_debug_frame_permission_frame_o2                   : out std_logic;
    fabric_debug_frame_permission_frame_o3                   : out std_logic;
    fabric_debug_frame_permission_frame_o4                   : out std_logic;
    fabric_otp_user_pwok_o                                   : out std_logic;
    fabric_otp_user_bend2_o                                  : out std_logic;
    fabric_mrepair_fuse_ded_o                                : out std_logic;
    fabric_debug_access_reg_data_ready_o                     : out std_logic;
    fabric_data_to_bist_o1                                   : out std_logic;
    fabric_data_to_bist_o2                                   : out std_logic;
    fabric_data_to_bist_o3                                   : out std_logic;
    fabric_data_to_bist_o4                                   : out std_logic;
    fabric_data_to_bist_o5                                   : out std_logic;
    fabric_data_to_bist_o6                                   : out std_logic;
    fabric_data_to_bist_o7                                   : out std_logic;
    fabric_data_to_bist_o8                                   : out std_logic;
    fabric_data_to_bist_o9                                   : out std_logic;
    fabric_data_to_bist_o10                                  : out std_logic;
    fabric_data_to_bist_o11                                  : out std_logic;
    fabric_data_to_bist_o12                                  : out std_logic;
    fabric_data_to_bist_o13                                  : out std_logic;
    fabric_data_to_bist_o14                                  : out std_logic;
    fabric_data_to_bist_o15                                  : out std_logic;
    fabric_data_to_bist_o16                                  : out std_logic;
    fabric_data_to_bist_o17                                  : out std_logic;
    fabric_data_to_bist_o18                                  : out std_logic;
    fabric_data_to_bist_o19                                  : out std_logic;
    fabric_data_to_bist_o20                                  : out std_logic;
    fabric_data_to_bist_o21                                  : out std_logic;
    fabric_data_to_bist_o22                                  : out std_logic;
    fabric_data_to_bist_o23                                  : out std_logic;
    fabric_data_to_bist_o24                                  : out std_logic;
    fabric_otp_user_startword_o1                             : out std_logic;
    fabric_otp_user_startword_o2                             : out std_logic;
    fabric_otp_user_startword_o3                             : out std_logic;
    fabric_otp_user_startword_o4                             : out std_logic;
    fabric_otp_user_startword_o5                             : out std_logic;
    fabric_otp_user_startword_o6                             : out std_logic;
    fabric_otp_user_startword_o7                             : out std_logic;
    fabric_otp_user_startword_o8                             : out std_logic;
    fabric_otp_user_startword_o9                             : out std_logic;
    fabric_otp_user_startword_o10                            : out std_logic;
    fabric_otp_user_startword_o11                            : out std_logic;
    fabric_otp_user_startword_o12                            : out std_logic;
    fabric_otp_user_startword_o13                            : out std_logic;
    fabric_otp_user_startword_o14                            : out std_logic;
    fabric_otp_user_startword_o15                            : out std_logic;
    fabric_otp_user_startword_o16                            : out std_logic;
    fabric_ahb_direct_data_o1                                : out std_logic;
    fabric_ahb_direct_data_o2                                : out std_logic;
    fabric_ahb_direct_data_o3                                : out std_logic;
    fabric_ahb_direct_data_o4                                : out std_logic;
    fabric_ahb_direct_data_o5                                : out std_logic;
    fabric_ahb_direct_data_o6                                : out std_logic;
    fabric_ahb_direct_data_o7                                : out std_logic;
    fabric_ahb_direct_data_o8                                : out std_logic;
    fabric_ahb_direct_data_o9                                : out std_logic;
    fabric_ahb_direct_data_o10                               : out std_logic;
    fabric_ahb_direct_data_o11                               : out std_logic;
    fabric_ahb_direct_data_o12                               : out std_logic;
    fabric_ahb_direct_data_o13                               : out std_logic;
    fabric_ahb_direct_data_o14                               : out std_logic;
    fabric_ahb_direct_data_o15                               : out std_logic;
    fabric_ahb_direct_data_o16                               : out std_logic;
    fabric_ahb_direct_data_o17                               : out std_logic;
    fabric_ahb_direct_data_o18                               : out std_logic;
    fabric_ahb_direct_data_o19                               : out std_logic;
    fabric_ahb_direct_data_o20                               : out std_logic;
    fabric_ahb_direct_data_o21                               : out std_logic;
    fabric_ahb_direct_data_o22                               : out std_logic;
    fabric_ahb_direct_data_o23                               : out std_logic;
    fabric_ahb_direct_data_o24                               : out std_logic;
    fabric_ahb_direct_data_o25                               : out std_logic;
    fabric_ahb_direct_data_o26                               : out std_logic;
    fabric_ahb_direct_data_o27                               : out std_logic;
    fabric_ahb_direct_data_o28                               : out std_logic;
    fabric_ahb_direct_data_o29                               : out std_logic;
    fabric_ahb_direct_data_o30                               : out std_logic;
    fabric_ahb_direct_data_o31                               : out std_logic;
    fabric_ahb_direct_data_o32                               : out std_logic;
    fabric_parusr_data_o1                                    : out std_logic;
    fabric_parusr_data_o2                                    : out std_logic;
    fabric_parusr_data_o3                                    : out std_logic;
    fabric_parusr_data_o4                                    : out std_logic;
    fabric_parusr_data_o5                                    : out std_logic;
    fabric_parusr_data_o6                                    : out std_logic;
    fabric_parusr_data_o7                                    : out std_logic;
    fabric_parusr_data_o8                                    : out std_logic;
    fabric_parusr_data_o9                                    : out std_logic;
    fabric_parusr_data_o10                                   : out std_logic;
    fabric_parusr_data_o11                                   : out std_logic;
    fabric_parusr_data_o12                                   : out std_logic;
    fabric_parusr_data_o13                                   : out std_logic;
    fabric_parusr_data_o14                                   : out std_logic;
    fabric_parusr_data_o15                                   : out std_logic;
    fabric_parusr_data_o16                                   : out std_logic;
    fabric_debug_otp_reload_err_o                            : out std_logic;
    fabric_cfg_fabric_user_unmask_o                          : out std_logic;
    fabric_decoder_init_ready_o                              : out std_logic;
    fabric_global_chip_status_o1                             : out std_logic;
    fabric_global_chip_status_o2                             : out std_logic;
    fabric_global_chip_status_o3                             : out std_logic;
    fabric_debug_security_boot_done_o                        : out std_logic;
    fabric_otp_user_calibrated_o                             : out std_logic;
    fabric_fuse_status_o1                                    : out std_logic;
    fabric_fuse_status_o2                                    : out std_logic;
    fabric_fuse_status_o3                                    : out std_logic;
    fabric_otp_apb_rdata_o1                                  : out std_logic;
    fabric_otp_apb_rdata_o2                                  : out std_logic;
    fabric_otp_apb_rdata_o3                                  : out std_logic;
    fabric_otp_apb_rdata_o4                                  : out std_logic;
    fabric_otp_apb_rdata_o5                                  : out std_logic;
    fabric_otp_apb_rdata_o6                                  : out std_logic;
    fabric_otp_apb_rdata_o7                                  : out std_logic;
    fabric_otp_apb_rdata_o8                                  : out std_logic;
    fabric_otp_apb_rdata_o9                                  : out std_logic;
    fabric_otp_apb_rdata_o10                                 : out std_logic;
    fabric_otp_apb_rdata_o11                                 : out std_logic;
    fabric_otp_apb_rdata_o12                                 : out std_logic;
    fabric_otp_apb_rdata_o13                                 : out std_logic;
    fabric_otp_apb_rdata_o14                                 : out std_logic;
    fabric_otp_apb_rdata_o15                                 : out std_logic;
    fabric_otp_apb_rdata_o16                                 : out std_logic;
    fabric_otp_apb_rdata_o17                                 : out std_logic;
    fabric_otp_apb_rdata_o18                                 : out std_logic;
    fabric_otp_apb_rdata_o19                                 : out std_logic;
    fabric_otp_apb_rdata_o20                                 : out std_logic;
    fabric_otp_apb_rdata_o21                                 : out std_logic;
    fabric_otp_apb_rdata_o22                                 : out std_logic;
    fabric_otp_apb_rdata_o23                                 : out std_logic;
    fabric_otp_apb_rdata_o24                                 : out std_logic;
    fabric_otp_apb_rdata_o25                                 : out std_logic;
    fabric_otp_apb_rdata_o26                                 : out std_logic;
    fabric_otp_apb_rdata_o27                                 : out std_logic;
    fabric_otp_apb_rdata_o28                                 : out std_logic;
    fabric_otp_apb_rdata_o29                                 : out std_logic;
    fabric_otp_apb_rdata_o30                                 : out std_logic;
    fabric_otp_apb_rdata_o31                                 : out std_logic;
    fabric_otp_apb_rdata_o32                                 : out std_logic;
    fabric_jtag_tms_o                                        : out std_logic;
    fabric_debug_bsec_core_status_o1                         : out std_logic;
    fabric_debug_bsec_core_status_o2                         : out std_logic;
    fabric_debug_bsec_core_status_o3                         : out std_logic;
    fabric_debug_bsec_core_status_o4                         : out std_logic;
    fabric_debug_bsec_core_status_o5                         : out std_logic;
    fabric_debug_bsec_core_status_o6                         : out std_logic;
    fabric_debug_bsec_core_status_o7                         : out std_logic;
    fabric_debug_bsec_core_status_o8                         : out std_logic;
    fabric_debug_bsec_core_status_o9                         : out std_logic;
    fabric_debug_bsec_core_status_o10                        : out std_logic;
    fabric_debug_bsec_core_status_o11                        : out std_logic;
    fabric_debug_bsec_core_status_o12                        : out std_logic;
    fabric_debug_bsec_core_status_o13                        : out std_logic;
    fabric_debug_bsec_core_status_o14                        : out std_logic;
    fabric_debug_bsec_core_status_o15                        : out std_logic;
    fabric_debug_bsec_core_status_o16                        : out std_logic;
    fabric_debug_bsec_core_status_o17                        : out std_logic;
    fabric_debug_bsec_core_status_o18                        : out std_logic;
    fabric_debug_bsec_core_status_o19                        : out std_logic;
    fabric_debug_bsec_core_status_o20                        : out std_logic;
    fabric_debug_bsec_core_status_o21                        : out std_logic;
    fabric_debug_bsec_core_status_o22                        : out std_logic;
    fabric_debug_bsec_core_status_o23                        : out std_logic;
    fabric_debug_bsec_core_status_o24                        : out std_logic;
    fabric_debug_bsec_core_status_o25                        : out std_logic;
    fabric_debug_bsec_core_status_o26                        : out std_logic;
    fabric_debug_bsec_core_status_o27                        : out std_logic;
    fabric_debug_bsec_core_status_o28                        : out std_logic;
    fabric_debug_bsec_core_status_o29                        : out std_logic;
    fabric_debug_bsec_core_status_o30                        : out std_logic;
    fabric_debug_bsec_core_status_o31                        : out std_logic;
    fabric_debug_bsec_core_status_o32                        : out std_logic;
    fabric_mrepair_fuse_bist1fail_o1                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o2                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o3                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o4                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o5                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o6                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o7                         : out std_logic;
    fabric_mrepair_fuse_bist1fail_o8                         : out std_logic;
    fabric_flag_ready_o                                      : out std_logic;
    fabric_mrepair_fuse_dout_o1                              : out std_logic;
    fabric_mrepair_fuse_dout_o2                              : out std_logic;
    fabric_mrepair_fuse_dout_o3                              : out std_logic;
    fabric_mrepair_fuse_dout_o4                              : out std_logic;
    fabric_mrepair_fuse_dout_o5                              : out std_logic;
    fabric_mrepair_fuse_dout_o6                              : out std_logic;
    fabric_mrepair_fuse_dout_o7                              : out std_logic;
    fabric_mrepair_fuse_dout_o8                              : out std_logic;
    fabric_mrepair_fuse_dout_o9                              : out std_logic;
    fabric_mrepair_fuse_dout_o10                             : out std_logic;
    fabric_mrepair_fuse_dout_o11                             : out std_logic;
    fabric_mrepair_fuse_dout_o12                             : out std_logic;
    fabric_mrepair_fuse_dout_o13                             : out std_logic;
    fabric_mrepair_fuse_dout_o14                             : out std_logic;
    fabric_mrepair_fuse_dout_o15                             : out std_logic;
    fabric_mrepair_fuse_dout_o16                             : out std_logic;
    fabric_mrepair_fuse_dout_o17                             : out std_logic;
    fabric_mrepair_fuse_dout_o18                             : out std_logic;
    fabric_mrepair_fuse_dout_o19                             : out std_logic;
    fabric_mrepair_fuse_dout_o20                             : out std_logic;
    fabric_mrepair_fuse_dout_o21                             : out std_logic;
    fabric_mrepair_fuse_dout_o22                             : out std_logic;
    fabric_mrepair_fuse_dout_o23                             : out std_logic;
    fabric_mrepair_fuse_dout_o24                             : out std_logic;
    fabric_mrepair_fuse_dout_o25                             : out std_logic;
    fabric_mrepair_fuse_dout_o26                             : out std_logic;
    fabric_mrepair_fuse_dout_o27                             : out std_logic;
    fabric_mrepair_fuse_dout_o28                             : out std_logic;
    fabric_mrepair_fuse_dout_o29                             : out std_logic;
    fabric_mrepair_fuse_dout_o30                             : out std_logic;
    fabric_mrepair_fuse_dout_o31                             : out std_logic;
    fabric_mrepair_fuse_dout_o32                             : out std_logic;
    fabric_mrepair_fuse_dout_o33                             : out std_logic;
    fabric_mrepair_fuse_dout_o34                             : out std_logic;
    fabric_mrepair_fuse_dout_o35                             : out std_logic;
    fabric_mrepair_fuse_dout_o36                             : out std_logic;
    fabric_mrepair_fuse_dout_o37                             : out std_logic;
    fabric_mrepair_fuse_dout_o38                             : out std_logic;
    fabric_mrepair_fuse_dout_o39                             : out std_logic;
    fabric_mrepair_fuse_dout_o40                             : out std_logic;
    fabric_mrepair_fuse_dout_o41                             : out std_logic;
    fabric_debug_rst_soft_o                                  : out std_logic;
    fabric_otp_user_ack_o                                    : out std_logic;
    fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o  : out std_logic;
    fabric_shift_en_to_bist_o1                               : out std_logic;
    fabric_shift_en_to_bist_o2                               : out std_logic;
    fabric_shift_en_to_bist_o3                               : out std_logic;
    fabric_shift_en_to_bist_o4                               : out std_logic;
    fabric_shift_en_to_bist_o5                               : out std_logic;
    fabric_shift_en_to_bist_o6                               : out std_logic;
    fabric_shift_en_to_bist_o7                               : out std_logic;
    fabric_shift_en_to_bist_o8                               : out std_logic;
    fabric_shift_en_to_bist_o9                               : out std_logic;
    fabric_shift_en_to_bist_o10                              : out std_logic;
    fabric_shift_en_to_bist_o11                              : out std_logic;
    fabric_shift_en_to_bist_o12                              : out std_logic;
    fabric_shift_en_to_bist_o13                              : out std_logic;
    fabric_shift_en_to_bist_o14                              : out std_logic;
    fabric_shift_en_to_bist_o15                              : out std_logic;
    fabric_shift_en_to_bist_o16                              : out std_logic;
    fabric_shift_en_to_bist_o17                              : out std_logic;
    fabric_shift_en_to_bist_o18                              : out std_logic;
    fabric_shift_en_to_bist_o19                              : out std_logic;
    fabric_shift_en_to_bist_o20                              : out std_logic;
    fabric_shift_en_to_bist_o21                              : out std_logic;
    fabric_shift_en_to_bist_o22                              : out std_logic;
    fabric_shift_en_to_bist_o23                              : out std_logic;
    fabric_shift_en_to_bist_o24                              : out std_logic;
    fabric_sif_reg_en_to_bist_o1                             : out std_logic;
    fabric_sif_reg_en_to_bist_o2                             : out std_logic;
    fabric_sif_reg_en_to_bist_o3                             : out std_logic;
    fabric_sif_reg_en_to_bist_o4                             : out std_logic;
    fabric_sif_reg_en_to_bist_o5                             : out std_logic;
    fabric_sif_reg_en_to_bist_o6                             : out std_logic;
    fabric_sif_reg_en_to_bist_o7                             : out std_logic;
    fabric_sif_reg_en_to_bist_o8                             : out std_logic;
    fabric_sif_reg_en_to_bist_o9                             : out std_logic;
    fabric_sif_reg_en_to_bist_o10                            : out std_logic;
    fabric_sif_reg_en_to_bist_o11                            : out std_logic;
    fabric_sif_reg_en_to_bist_o12                            : out std_logic;
    fabric_sif_reg_en_to_bist_o13                            : out std_logic;
    fabric_sif_reg_en_to_bist_o14                            : out std_logic;
    fabric_sif_reg_en_to_bist_o15                            : out std_logic;
    fabric_sif_reg_en_to_bist_o16                            : out std_logic;
    fabric_sif_reg_en_to_bist_o17                            : out std_logic;
    fabric_sif_reg_en_to_bist_o18                            : out std_logic;
    fabric_sif_reg_en_to_bist_o19                            : out std_logic;
    fabric_sif_reg_en_to_bist_o20                            : out std_logic;
    fabric_sif_reg_en_to_bist_o21                            : out std_logic;
    fabric_sif_reg_en_to_bist_o22                            : out std_logic;
    fabric_sif_reg_en_to_bist_o23                            : out std_logic;
    fabric_sif_reg_en_to_bist_o24                            : out std_logic;
    fabric_sif_reg_en_to_bist_o25                            : out std_logic;
    fabric_sif_reg_en_to_bist_o26                            : out std_logic;
    fabric_sif_reg_en_to_bist_o27                            : out std_logic;
    fabric_sif_reg_en_to_bist_o28                            : out std_logic;
    fabric_sif_reg_en_to_bist_o29                            : out std_logic;
    fabric_sif_reg_en_to_bist_o30                            : out std_logic;
    fabric_sif_reg_en_to_bist_o31                            : out std_logic;
    fabric_sif_reg_en_to_bist_o32                            : out std_logic;
    fabric_sif_reg_en_to_bist_o33                            : out std_logic;
    fabric_sif_reg_en_to_bist_o34                            : out std_logic;
    fabric_sif_reg_en_to_bist_o35                            : out std_logic;
    fabric_sif_reg_en_to_bist_o36                            : out std_logic;
    fabric_sif_reg_en_to_bist_o37                            : out std_logic;
    fabric_sif_reg_en_to_bist_o38                            : out std_logic;
    fabric_sif_reg_en_to_bist_o39                            : out std_logic;
    fabric_sif_reg_en_to_bist_o40                            : out std_logic;
    fabric_sif_reg_en_to_bist_o41                            : out std_logic;
    fabric_sif_reg_en_to_bist_o42                            : out std_logic;
    fabric_sif_reg_en_to_bist_o43                            : out std_logic;
    fabric_sif_reg_en_to_bist_o44                            : out std_logic;
    fabric_sif_reg_en_to_bist_o45                            : out std_logic;
    fabric_sif_reg_en_to_bist_o46                            : out std_logic;
    fabric_sif_reg_en_to_bist_o47                            : out std_logic;
    fabric_sif_reg_en_to_bist_o48                            : out std_logic;
    fabric_sif_reg_en_to_bist_o49                            : out std_logic;
    fabric_sif_reg_en_to_bist_o50                            : out std_logic;
    fabric_sif_reg_en_to_bist_o51                            : out std_logic;
    fabric_sif_reg_en_to_bist_o52                            : out std_logic;
    fabric_sif_reg_en_to_bist_o53                            : out std_logic;
    fabric_sif_reg_en_to_bist_o54                            : out std_logic;
    fabric_sif_reg_en_to_bist_o55                            : out std_logic;
    fabric_sif_reg_en_to_bist_o56                            : out std_logic;
    fabric_sif_reg_en_to_bist_o57                            : out std_logic;
    fabric_sif_reg_en_to_bist_o58                            : out std_logic;
    fabric_sif_reg_en_to_bist_o59                            : out std_logic;
    fabric_sif_reg_en_to_bist_o60                            : out std_logic;
    fabric_sif_reg_en_to_bist_o61                            : out std_logic;
    fabric_sif_reg_en_to_bist_o62                            : out std_logic;
    fabric_sif_reg_en_to_bist_o63                            : out std_logic;
    fabric_sif_reg_en_to_bist_o64                            : out std_logic;
    fabric_sif_reg_en_to_bist_o65                            : out std_logic;
    fabric_sif_reg_en_to_bist_o66                            : out std_logic;
    fabric_sif_reg_en_to_bist_o67                            : out std_logic;
    fabric_sif_reg_en_to_bist_o68                            : out std_logic;
    fabric_sif_reg_en_to_bist_o69                            : out std_logic;
    fabric_sif_reg_en_to_bist_o70                            : out std_logic;
    fabric_sif_reg_en_to_bist_o71                            : out std_logic;
    fabric_sif_reg_en_to_bist_o72                            : out std_logic;
    fabric_sif_reg_en_to_bist_o73                            : out std_logic;
    fabric_sif_reg_en_to_bist_o74                            : out std_logic;
    fabric_sif_reg_en_to_bist_o75                            : out std_logic;
    fabric_sif_reg_en_to_bist_o76                            : out std_logic;
    fabric_sif_reg_en_to_bist_o77                            : out std_logic;
    fabric_sif_reg_en_to_bist_o78                            : out std_logic;
    fabric_sif_reg_en_to_bist_o79                            : out std_logic;
    fabric_sif_reg_en_to_bist_o80                            : out std_logic;
    fabric_sif_reg_en_to_bist_o81                            : out std_logic;
    fabric_sif_reg_en_to_bist_o82                            : out std_logic;
    fabric_sif_reg_en_to_bist_o83                            : out std_logic;
    fabric_sif_reg_en_to_bist_o84                            : out std_logic;
    fabric_sif_reg_en_to_bist_o85                            : out std_logic;
    fabric_sif_reg_en_to_bist_o86                            : out std_logic;
    fabric_sif_reg_en_to_bist_o87                            : out std_logic;
    fabric_sif_reg_en_to_bist_o88                            : out std_logic;
    fabric_sif_reg_en_to_bist_o89                            : out std_logic;
    fabric_sif_reg_en_to_bist_o90                            : out std_logic;
    fabric_sif_reg_en_to_bist_o91                            : out std_logic;
    fabric_sif_reg_en_to_bist_o92                            : out std_logic;
    fabric_sif_reg_en_to_bist_o93                            : out std_logic;
    fabric_sif_reg_en_to_bist_o94                            : out std_logic;
    fabric_sif_reg_en_to_bist_o95                            : out std_logic;
    fabric_sif_reg_en_to_bist_o96                            : out std_logic;
    fabric_sif_reg_en_to_bist_o97                            : out std_logic;
    fabric_sif_reg_en_to_bist_o98                            : out std_logic;
    fabric_sif_reg_en_to_bist_o99                            : out std_logic;
    fabric_sif_reg_en_to_bist_o100                           : out std_logic;
    fabric_sif_reg_en_to_bist_o101                           : out std_logic;
    fabric_sif_reg_en_to_bist_o102                           : out std_logic;
    fabric_sif_reg_en_to_bist_o103                           : out std_logic;
    fabric_sif_reg_en_to_bist_o104                           : out std_logic;
    fabric_sif_reg_en_to_bist_o105                           : out std_logic;
    fabric_sif_reg_en_to_bist_o106                           : out std_logic;
    fabric_sif_reg_en_to_bist_o107                           : out std_logic;
    fabric_sif_reg_en_to_bist_o108                           : out std_logic;
    fabric_sif_reg_en_to_bist_o109                           : out std_logic;
    fabric_sif_reg_en_to_bist_o110                           : out std_logic;
    fabric_sif_reg_en_to_bist_o111                           : out std_logic;
    fabric_sif_reg_en_to_bist_o112                           : out std_logic;
    fabric_sif_reg_en_to_bist_o113                           : out std_logic;
    fabric_sif_reg_en_to_bist_o114                           : out std_logic;
    fabric_sif_reg_en_to_bist_o115                           : out std_logic;
    fabric_sif_reg_en_to_bist_o116                           : out std_logic;
    fabric_sif_reg_en_to_bist_o117                           : out std_logic;
    fabric_sif_reg_en_to_bist_o118                           : out std_logic;
    fabric_sif_reg_en_to_bist_o119                           : out std_logic;
    fabric_sif_reg_en_to_bist_o120                           : out std_logic;
    fabric_debug_otp_manager_read_otp_o                      : out std_logic;
    fabric_otp_user_sec_o                                    : out std_logic;
    fabric_otp_user_wlromout_o1                              : out std_logic;
    fabric_otp_user_wlromout_o2                              : out std_logic;
    fabric_otp_user_wlromout_o3                              : out std_logic;
    fabric_otp_user_wlromout_o4                              : out std_logic;
    fabric_otp_user_wlromout_o5                              : out std_logic;
    fabric_otp_user_wlromout_o6                              : out std_logic;
    fabric_otp_user_wlromout_o7                              : out std_logic;
    fabric_otp_user_wlromout_o8                              : out std_logic;
    fabric_otp_user_wlromout_o9                              : out std_logic;
    fabric_otp_user_wlromout_o10                             : out std_logic;
    fabric_mrepair_fuse_bend1_o                              : out std_logic;
    fabric_mrepair_fuse_flagstate_o1                         : out std_logic;
    fabric_mrepair_fuse_flagstate_o2                         : out std_logic;
    fabric_mrepair_fuse_flagstate_o3                         : out std_logic;
    fabric_mrepair_fuse_flagstate_o4                         : out std_logic;
    fabric_system_data_from_mem_bist_o1                      : out std_logic;
    fabric_system_data_from_mem_bist_o2                      : out std_logic;
    fabric_system_data_from_mem_bist_o3                      : out std_logic;
    fabric_system_data_from_mem_bist_o4                      : out std_logic;
    fabric_system_data_from_mem_bist_o5                      : out std_logic;
    fabric_system_data_from_mem_bist_o6                      : out std_logic;
    fabric_system_data_from_mem_bist_o7                      : out std_logic;
    fabric_system_data_from_mem_bist_o8                      : out std_logic;
    fabric_system_data_from_mem_bist_o9                      : out std_logic;
    fabric_system_data_from_mem_bist_o10                     : out std_logic;
    fabric_system_data_from_mem_bist_o11                     : out std_logic;
    fabric_system_data_from_mem_bist_o12                     : out std_logic;
    fabric_system_data_from_mem_bist_o13                     : out std_logic;
    fabric_system_data_from_mem_bist_o14                     : out std_logic;
    fabric_system_data_from_mem_bist_o15                     : out std_logic;
    fabric_system_data_from_mem_bist_o16                     : out std_logic;
    fabric_system_data_from_mem_bist_o17                     : out std_logic;
    fabric_system_data_from_mem_bist_o18                     : out std_logic;
    fabric_system_data_from_mem_bist_o19                     : out std_logic;
    fabric_system_data_from_mem_bist_o20                     : out std_logic;
    fabric_system_data_from_mem_bist_o21                     : out std_logic;
    fabric_system_data_from_mem_bist_o22                     : out std_logic;
    fabric_system_data_from_mem_bist_o23                     : out std_logic;
    fabric_system_data_from_mem_bist_o24                     : out std_logic;
    fabric_direct_data_o1                                    : out std_logic;
    fabric_direct_data_o2                                    : out std_logic;
    fabric_direct_data_o3                                    : out std_logic;
    fabric_direct_data_o4                                    : out std_logic;
    fabric_direct_data_o5                                    : out std_logic;
    fabric_direct_data_o6                                    : out std_logic;
    fabric_direct_data_o7                                    : out std_logic;
    fabric_direct_data_o8                                    : out std_logic;
    fabric_direct_data_o9                                    : out std_logic;
    fabric_direct_data_o10                                   : out std_logic;
    fabric_direct_data_o11                                   : out std_logic;
    fabric_direct_data_o12                                   : out std_logic;
    fabric_direct_data_o13                                   : out std_logic;
    fabric_direct_data_o14                                   : out std_logic;
    fabric_direct_data_o15                                   : out std_logic;
    fabric_direct_data_o16                                   : out std_logic;
    fabric_direct_data_o17                                   : out std_logic;
    fabric_direct_data_o18                                   : out std_logic;
    fabric_direct_data_o19                                   : out std_logic;
    fabric_direct_data_o20                                   : out std_logic;
    fabric_direct_data_o21                                   : out std_logic;
    fabric_direct_data_o22                                   : out std_logic;
    fabric_direct_data_o23                                   : out std_logic;
    fabric_direct_data_o24                                   : out std_logic;
    fabric_direct_data_o25                                   : out std_logic;
    fabric_direct_data_o26                                   : out std_logic;
    fabric_direct_data_o27                                   : out std_logic;
    fabric_direct_data_o28                                   : out std_logic;
    fabric_direct_data_o29                                   : out std_logic;
    fabric_direct_data_o30                                   : out std_logic;
    fabric_direct_data_o31                                   : out std_logic;
    fabric_direct_data_o32                                   : out std_logic;
    fabric_otp_user_bbad_o                                   : out std_logic;
    fabric_user_read_cycle_o                                 : out std_logic;
    fabric_chip_status_o1                                    : out std_logic;
    fabric_chip_status_o2                                    : out std_logic;
    fabric_chip_status_o3                                    : out std_logic;
    fabric_chip_status_o4                                    : out std_logic;
    fabric_chip_status_o5                                    : out std_logic;
    fabric_chip_status_o6                                    : out std_logic;
    fabric_chip_status_o7                                    : out std_logic;
    fabric_chip_status_o8                                    : out std_logic;
    fabric_chip_status_o9                                    : out std_logic;
    fabric_chip_status_o10                                   : out std_logic;
    fabric_chip_status_o11                                   : out std_logic;
    fabric_chip_status_o12                                   : out std_logic;
    fabric_chip_status_o13                                   : out std_logic;
    fabric_chip_status_o14                                   : out std_logic;
    fabric_chip_status_o15                                   : out std_logic;
    fabric_chip_status_o16                                   : out std_logic;
    fabric_chip_status_o17                                   : out std_logic;
    fabric_chip_status_o18                                   : out std_logic;
    fabric_chip_status_o19                                   : out std_logic;
    fabric_chip_status_o20                                   : out std_logic;
    fabric_chip_status_o21                                   : out std_logic;
    fabric_chip_status_o22                                   : out std_logic;
    fabric_chip_status_o23                                   : out std_logic;
    fabric_chip_status_o24                                   : out std_logic;
    fabric_chip_status_o25                                   : out std_logic;
    fabric_chip_status_o26                                   : out std_logic;
    fabric_chip_status_o27                                   : out std_logic;
    fabric_chip_status_o28                                   : out std_logic;
    fabric_chip_status_o29                                   : out std_logic;
    fabric_chip_status_o30                                   : out std_logic;
    fabric_chip_status_o31                                   : out std_logic;
    fabric_chip_status_o32                                   : out std_logic;
    fabric_chip_status_o33                                   : out std_logic;
    fabric_chip_status_o34                                   : out std_logic;
    fabric_chip_status_o35                                   : out std_logic;
    fabric_chip_status_o36                                   : out std_logic;
    fabric_chip_status_o37                                   : out std_logic;
    fabric_chip_status_o38                                   : out std_logic;
    fabric_chip_status_o39                                   : out std_logic;
    fabric_chip_status_o40                                   : out std_logic;
    fabric_chip_status_o41                                   : out std_logic;
    fabric_chip_status_o42                                   : out std_logic;
    fabric_chip_status_o43                                   : out std_logic;
    fabric_chip_status_o44                                   : out std_logic;
    fabric_chip_status_o45                                   : out std_logic;
    fabric_chip_status_o46                                   : out std_logic;
    fabric_chip_status_o47                                   : out std_logic;
    fabric_chip_status_o48                                   : out std_logic;
    fabric_chip_status_o49                                   : out std_logic;
    fabric_chip_status_o50                                   : out std_logic;
    fabric_chip_status_o51                                   : out std_logic;
    fabric_chip_status_o52                                   : out std_logic;
    fabric_chip_status_o53                                   : out std_logic;
    fabric_chip_status_o54                                   : out std_logic;
    fabric_chip_status_o55                                   : out std_logic;
    fabric_chip_status_o56                                   : out std_logic;
    fabric_chip_status_o57                                   : out std_logic;
    fabric_chip_status_o58                                   : out std_logic;
    fabric_chip_status_o59                                   : out std_logic;
    fabric_chip_status_o60                                   : out std_logic;
    fabric_chip_status_o61                                   : out std_logic;
    fabric_chip_status_o62                                   : out std_logic;
    fabric_chip_status_o63                                   : out std_logic;
    fabric_chip_status_o64                                   : out std_logic;
    fabric_chip_status_o65                                   : out std_logic;
    fabric_chip_status_o66                                   : out std_logic;
    fabric_chip_status_o67                                   : out std_logic;
    fabric_chip_status_o68                                   : out std_logic;
    fabric_chip_status_o69                                   : out std_logic;
    fabric_chip_status_o70                                   : out std_logic;
    fabric_chip_status_o71                                   : out std_logic;
    fabric_chip_status_o72                                   : out std_logic;
    fabric_mrepair_fuse_disturbed_o                          : out std_logic;
    fabric_debug_otpboot_state_o1                            : out std_logic;
    fabric_debug_otpboot_state_o2                            : out std_logic;
    fabric_debug_otpboot_state_o3                            : out std_logic;
    fabric_pd_ready_o1                                       : out std_logic;
    fabric_pd_ready_o2                                       : out std_logic;
    fabric_pd_ready_o3                                       : out std_logic;
    fabric_pd_ready_o4                                       : out std_logic;
    fabric_pd_ready_o5                                       : out std_logic;
    fabric_pd_ready_o6                                       : out std_logic;
    fabric_pd_ready_o7                                       : out std_logic;
    fabric_pd_ready_o8                                       : out std_logic;
    fabric_pd_ready_o9                                       : out std_logic;
    fabric_pd_ready_o10                                      : out std_logic;
    fabric_pd_ready_o11                                      : out std_logic;
    fabric_pd_ready_o12                                      : out std_logic;
    fabric_pd_ready_o13                                      : out std_logic;
    fabric_pd_ready_o14                                      : out std_logic;
    fabric_pd_ready_o15                                      : out std_logic;
    fabric_pd_ready_o16                                      : out std_logic;
    fabric_pd_ready_o17                                      : out std_logic;
    fabric_pd_ready_o18                                      : out std_logic;
    fabric_pd_ready_o19                                      : out std_logic;
    fabric_pd_ready_o20                                      : out std_logic;
    fabric_pd_ready_o21                                      : out std_logic;
    fabric_pd_ready_o22                                      : out std_logic;
    fabric_pd_ready_o23                                      : out std_logic;
    fabric_pd_ready_o24                                      : out std_logic;
    fabric_debug_key_correct_o                               : out std_logic;
    fabric_otp_apb_ready_o                                   : out std_logic;
    fabric_otp_user_progfail_o                               : out std_logic;
    fabric_mrepair_fuse_sec_o                                : out std_logic;
    fabric_mrepair_fuse_bend2_o                              : out std_logic;
    fabric_debug_lifecycle_o1                                : out std_logic;
    fabric_debug_lifecycle_o2                                : out std_logic;
    fabric_debug_lifecycle_o3                                : out std_logic;
    fabric_debug_lifecycle_o4                                : out std_logic;
    fabric_mrepair_fuse_ack_o                                : out std_logic;
    fabric_debug_cpt_retry_o1                                : out std_logic;
    fabric_debug_cpt_retry_o2                                : out std_logic;
    fabric_debug_cpt_retry_o3                                : out std_logic;
    fabric_debug_cpt_retry_o4                                : out std_logic;
    fabric_otp_security_ack_o                                : out std_logic;
    fabric_debug_otpmgmt_state_o1                            : out std_logic;
    fabric_debug_otpmgmt_state_o2                            : out std_logic;
    fabric_debug_otpmgmt_state_o3                            : out std_logic;
    fabric_mrepair_fuse_progfail_o                           : out std_logic;
    fabric_otp_user_bist2fail_o1                             : out std_logic;
    fabric_otp_user_bist2fail_o2                             : out std_logic;
    fabric_otp_user_bist2fail_o3                             : out std_logic;
    fabric_otp_user_bist2fail_o4                             : out std_logic;
    fabric_otp_user_bist2fail_o5                             : out std_logic;
    fabric_otp_user_bist2fail_o6                             : out std_logic;
    fabric_otp_user_bist2fail_o7                             : out std_logic;
    fabric_user_data_o1                                      : out std_logic;
    fabric_user_data_o2                                      : out std_logic;
    fabric_user_data_o3                                      : out std_logic;
    fabric_user_data_o4                                      : out std_logic;
    fabric_user_data_o5                                      : out std_logic;
    fabric_user_data_o6                                      : out std_logic;
    fabric_user_data_o7                                      : out std_logic;
    fabric_user_data_o8                                      : out std_logic;
    fabric_user_data_o9                                      : out std_logic;
    fabric_user_data_o10                                     : out std_logic;
    fabric_user_data_o11                                     : out std_logic;
    fabric_user_data_o12                                     : out std_logic;
    fabric_user_data_o13                                     : out std_logic;
    fabric_user_data_o14                                     : out std_logic;
    fabric_user_data_o15                                     : out std_logic;
    fabric_user_data_o16                                     : out std_logic;
    fabric_user_data_o17                                     : out std_logic;
    fabric_user_data_o18                                     : out std_logic;
    fabric_user_data_o19                                     : out std_logic;
    fabric_user_data_o20                                     : out std_logic;
    fabric_user_data_o21                                     : out std_logic;
    fabric_user_data_o22                                     : out std_logic;
    fabric_user_data_o23                                     : out std_logic;
    fabric_user_data_o24                                     : out std_logic;
    fabric_user_data_o25                                     : out std_logic;
    fabric_user_data_o26                                     : out std_logic;
    fabric_user_data_o27                                     : out std_logic;
    fabric_user_data_o28                                     : out std_logic;
    fabric_user_data_o29                                     : out std_logic;
    fabric_user_data_o30                                     : out std_logic;
    fabric_user_data_o31                                     : out std_logic;
    fabric_user_data_o32                                     : out std_logic;
    fabric_jtag_tdi_o                                        : out std_logic;
    fabric_lowskew_o3                                        : out std_logic;
    fabric_lowskew_o5                                        : out std_logic;
    fabric_lowskew_o4                                        : out std_logic;
    fabric_debug_error_o                                     : out std_logic;
    fabric_jtag_usr2_o                                       : out std_logic;
    fabric_mrepair_fuse_wlromout_o1                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o2                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o3                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o4                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o5                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o6                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o7                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o8                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o9                          : out std_logic;
    fabric_mrepair_fuse_wlromout_o10                         : out std_logic;
    fabric_debug_otpapb_state_o1                             : out std_logic;
    fabric_debug_otpapb_state_o2                             : out std_logic;
    fabric_debug_otpapb_state_o3                             : out std_logic;
    fabric_otp_user_bist1fail_o1                             : out std_logic;
    fabric_otp_user_bist1fail_o2                             : out std_logic;
    fabric_otp_user_bist1fail_o3                             : out std_logic;
    fabric_otp_user_bist1fail_o4                             : out std_logic;
    fabric_otp_user_bist1fail_o5                             : out std_logic;
    fabric_otp_user_bist1fail_o6                             : out std_logic;
    fabric_otp_user_bist1fail_o7                             : out std_logic;
    fabric_otp_user_bist1fail_o8                             : out std_logic;
    fabric_otp_security_bist_fail2_o1                        : out std_logic;
    fabric_otp_security_bist_fail2_o2                        : out std_logic;
    fabric_otp_security_bist_fail2_o3                        : out std_logic;
    fabric_otp_security_bist_fail2_o4                        : out std_logic;
    fabric_otp_security_bist_fail2_o5                        : out std_logic;
    fabric_otp_security_bist_fail2_o6                        : out std_logic;
    fabric_otp_security_bist_fail2_o7                        : out std_logic;
    fabric_otp_user_disturbed_o                              : out std_logic;
    fabric_flag_trigger_o                                    : out std_logic;
    fabric_otp_security_bist_end2_o                          : out std_logic;
    fabric_otp_security_bist_fail1_o1                        : out std_logic;
    fabric_otp_security_bist_fail1_o2                        : out std_logic;
    fabric_otp_security_bist_fail1_o3                        : out std_logic;
    fabric_otp_security_bist_fail1_o4                        : out std_logic;
    fabric_otp_security_bist_fail1_o5                        : out std_logic;
    fabric_otp_security_bist_fail1_o6                        : out std_logic;
    fabric_otp_security_bist_fail1_o7                        : out std_logic;
    fabric_otp_security_bist_fail1_o8                        : out std_logic;
    fabric_mrepair_fuse_locked_o                             : out std_logic;
    fabric_otp_user_flagstate_o1                             : out std_logic;
    fabric_otp_user_flagstate_o2                             : out std_logic;
    fabric_otp_user_flagstate_o3                             : out std_logic;
    fabric_otp_user_flagstate_o4                             : out std_logic;
    fabric_otp_security_scanout_o1                           : out std_logic;
    fabric_otp_security_scanout_o2                           : out std_logic;
    fabric_otp_security_scanout_o3                           : out std_logic;
    fabric_otp_security_scanout_o4                           : out std_logic;
    fabric_otp_security_scanout_o5                           : out std_logic;
    fabric_user_write_cycle_o                                : out std_logic;
    fabric_debug_fsm_state_o1                                : out std_logic;
    fabric_debug_fsm_state_o2                                : out std_logic;
    fabric_debug_fsm_state_o3                                : out std_logic;
    fabric_otp_user_ded_o                                    : out std_logic;
    fabric_debug_otp_manager_read_done_o                     : out std_logic;
    fabric_debug_frame_use_encryption_o                      : out std_logic;
    fabric_data_to_system_o                                  : out std_logic;
    fabric_jtag_usr1_o                                       : out std_logic;
    fabric_otp_user_bend1_o                                  : out std_logic;
    fabric_debug_otpboot_curr_addr_o1                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o2                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o3                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o4                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o5                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o6                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o7                        : out std_logic;
    fabric_debug_otpboot_curr_addr_o8                        : out std_logic;
    fabric_mrepair_fuse_ready_o                              : out std_logic;
    fabric_mrepair_fuse_calibrated_o                         : out std_logic;
    fabric_sif_load_en_to_bist_o1                            : out std_logic;
    fabric_sif_load_en_to_bist_o2                            : out std_logic;
    fabric_sif_load_en_to_bist_o3                            : out std_logic;
    fabric_sif_load_en_to_bist_o4                            : out std_logic;
    fabric_sif_load_en_to_bist_o5                            : out std_logic;
    fabric_sif_load_en_to_bist_o6                            : out std_logic;
    fabric_sif_load_en_to_bist_o7                            : out std_logic;
    fabric_sif_load_en_to_bist_o8                            : out std_logic;
    fabric_sif_load_en_to_bist_o9                            : out std_logic;
    fabric_sif_load_en_to_bist_o10                           : out std_logic;
    fabric_sif_load_en_to_bist_o11                           : out std_logic;
    fabric_sif_load_en_to_bist_o12                           : out std_logic;
    fabric_sif_load_en_to_bist_o13                           : out std_logic;
    fabric_sif_load_en_to_bist_o14                           : out std_logic;
    fabric_sif_load_en_to_bist_o15                           : out std_logic;
    fabric_sif_load_en_to_bist_o16                           : out std_logic;
    fabric_sif_load_en_to_bist_o17                           : out std_logic;
    fabric_sif_load_en_to_bist_o18                           : out std_logic;
    fabric_sif_load_en_to_bist_o19                           : out std_logic;
    fabric_sif_load_en_to_bist_o20                           : out std_logic;
    fabric_sif_load_en_to_bist_o21                           : out std_logic;
    fabric_sif_load_en_to_bist_o22                           : out std_logic;
    fabric_sif_load_en_to_bist_o23                           : out std_logic;
    fabric_sif_load_en_to_bist_o24                           : out std_logic;
    fabric_io_out_o1                                         : out std_logic;
    fabric_io_out_o2                                         : out std_logic;
    fabric_io_out_o3                                         : out std_logic;
    fabric_io_out_o4                                         : out std_logic;
    fabric_io_out_o5                                         : out std_logic;
    fabric_io_out_o6                                         : out std_logic;
    fabric_io_out_o7                                         : out std_logic;
    fabric_io_out_o8                                         : out std_logic;
    fabric_io_out_o9                                         : out std_logic;
    fabric_io_out_o10                                        : out std_logic;
    fabric_io_out_o11                                        : out std_logic;
    fabric_io_out_o12                                        : out std_logic;
    fabric_io_out_o13                                        : out std_logic;
    fabric_io_out_o14                                        : out std_logic;
    fabric_io_out_o15                                        : out std_logic;
    fabric_io_out_o16                                        : out std_logic;
    fabric_io_out_o17                                        : out std_logic;
    fabric_io_out_o18                                        : out std_logic;
    fabric_io_out_o19                                        : out std_logic;
    fabric_io_out_o20                                        : out std_logic;
    fabric_io_out_o21                                        : out std_logic;
    fabric_io_out_o22                                        : out std_logic;
    fabric_io_out_o23                                        : out std_logic;
    fabric_io_out_o24                                        : out std_logic;
    fabric_io_out_o25                                        : out std_logic;
    fabric_mrepair_fuse_startword_o1                         : out std_logic;
    fabric_mrepair_fuse_startword_o2                         : out std_logic;
    fabric_mrepair_fuse_startword_o3                         : out std_logic;
    fabric_mrepair_fuse_startword_o4                         : out std_logic;
    fabric_mrepair_fuse_startword_o5                         : out std_logic;
    fabric_mrepair_fuse_startword_o6                         : out std_logic;
    fabric_mrepair_fuse_startword_o7                         : out std_logic;
    fabric_mrepair_fuse_startword_o8                         : out std_logic;
    fabric_mrepair_fuse_startword_o9                         : out std_logic;
    fabric_mrepair_fuse_startword_o10                        : out std_logic;
    fabric_mrepair_fuse_startword_o11                        : out std_logic;
    fabric_mrepair_fuse_startword_o12                        : out std_logic;
    fabric_mrepair_fuse_startword_o13                        : out std_logic;
    fabric_mrepair_fuse_startword_o14                        : out std_logic;
    fabric_mrepair_fuse_startword_o15                        : out std_logic;
    fabric_mrepair_fuse_startword_o16                        : out std_logic;
    fabric_system_dataready_o                                : out std_logic;
    fabric_mrepair_fuse_pwok_o                               : out std_logic;
    fabric_lowskew_o6                                        : out std_logic;
    fabric_cfg_fabric_user_flag_o                            : out std_logic;
    fabric_otp_user_dout_o1                                  : out std_logic;
    fabric_otp_user_dout_o2                                  : out std_logic;
    fabric_otp_user_dout_o3                                  : out std_logic;
    fabric_otp_user_dout_o4                                  : out std_logic;
    fabric_otp_user_dout_o5                                  : out std_logic;
    fabric_otp_user_dout_o6                                  : out std_logic;
    fabric_otp_user_dout_o7                                  : out std_logic;
    fabric_otp_user_dout_o8                                  : out std_logic;
    fabric_otp_user_dout_o9                                  : out std_logic;
    fabric_otp_user_dout_o10                                 : out std_logic;
    fabric_otp_user_dout_o11                                 : out std_logic;
    fabric_otp_user_dout_o12                                 : out std_logic;
    fabric_otp_user_dout_o13                                 : out std_logic;
    fabric_otp_user_dout_o14                                 : out std_logic;
    fabric_otp_user_dout_o15                                 : out std_logic;
    fabric_otp_user_dout_o16                                 : out std_logic;
    fabric_otp_user_dout_o17                                 : out std_logic;
    fabric_otp_user_dout_o18                                 : out std_logic;
    fabric_otp_user_dout_o19                                 : out std_logic;
    fabric_otp_user_dout_o20                                 : out std_logic;
    fabric_otp_user_dout_o21                                 : out std_logic;
    fabric_otp_user_dout_o22                                 : out std_logic;
    fabric_otp_user_dout_o23                                 : out std_logic;
    fabric_otp_user_dout_o24                                 : out std_logic;
    fabric_otp_user_dout_o25                                 : out std_logic;
    fabric_otp_user_dout_o26                                 : out std_logic;
    fabric_otp_user_dout_o27                                 : out std_logic;
    fabric_otp_user_dout_o28                                 : out std_logic;
    fabric_otp_user_dout_o29                                 : out std_logic;
    fabric_otp_user_dout_o30                                 : out std_logic;
    fabric_otp_user_dout_o31                                 : out std_logic;
    fabric_otp_user_dout_o32                                 : out std_logic;
    fabric_otp_user_dout_o33                                 : out std_logic;
    fabric_otp_user_dout_o34                                 : out std_logic;
    fabric_otp_user_dout_o35                                 : out std_logic;
    fabric_otp_user_dout_o36                                 : out std_logic;
    fabric_otp_user_dout_o37                                 : out std_logic;
    fabric_otp_user_dout_o38                                 : out std_logic;
    fabric_otp_user_dout_o39                                 : out std_logic;
    fabric_otp_user_dout_o40                                 : out std_logic;
    fabric_otp_user_dout_o41                                 : out std_logic;
    fabric_mrepair_fuse_bist2fail_o1                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o2                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o3                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o4                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o5                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o6                         : out std_logic;
    fabric_mrepair_fuse_bist2fail_o7                         : out std_logic;
    fabric_status_cold_start_o                               : out std_logic;
    fabric_flag_error_o                                      : out std_logic;
    fabric_debug_direct_permission_read_o1                   : out std_logic;
    fabric_debug_direct_permission_read_o2                   : out std_logic;
    fabric_debug_direct_permission_read_o3                   : out std_logic;
    fabric_debug_direct_permission_read_o4                   : out std_logic
);
end NX_SERVICE_U;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--  NX_SERVICE_U_WRAP definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library NX;
use NX.nxPackage.all;
entity NX_SERVICE_U_WRAP is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    fabric_otp_user_tst_scanenable_i                         : in std_logic;
    fabric_otp_cfg_loader_read_en_i                          : in std_logic;
    fabric_otp_security_force_pdn1_i                         : in std_logic;
    fabric_otp_security_scanenable_i                         : in std_logic;
    fabric_otp_user_din_i                                    : in std_logic_vector(38 downto 0);
    fabric_mrepair_fuse_prgwidth_i                           : in std_logic_vector(2 downto 0);
    fabric_otp_apb_wdata_i                                   : in std_logic_vector(31 downto 0);
    fabric_otp_cfg_clk_otpm_disable_i                        : in std_logic;
    fabric_otp_user_disturbcheck_i                           : in std_logic;
    fabric_mrepair_fuse_read_i                               : in std_logic;
    fabric_otp_user_rbact2_i                                 : in std_logic;
    fabric_mrepair_fuse_eccbypass_i                          : in std_logic;
    fabric_otp_user_bistmode_i                               : in std_logic;
    fabric_otp_user_add_i                                    : in std_logic_vector(6 downto 0);
    fabric_otp_user_tm_i                                     : in std_logic;
    fabric_otp_rstn_i                                        : in std_logic;
    fabric_mrepair_fuse_disturbchecked_i                     : in std_logic;
    fabric_otp_user_rbact1_i                                 : in std_logic;
    fabric_mrepair_fuse_tst_scanin_i                         : in std_logic_vector(4 downto 0);
    fabric_parusr_type_i                                     : in std_logic_vector(1 downto 0);
    fabric_mrepair_fuse_redbypass_i                          : in std_logic;
    fabric_otp_user_eccbypass_i                              : in std_logic;
    fabric_otp_user_redbypass_i                              : in std_logic;
    fabric_mrepair_mode_i                                    : in std_logic_vector(3 downto 0);
    fabric_parusr_cs_i                                       : in std_logic;
    fabric_sif_reg_en_i                                      : in std_logic_vector(119 downto 0);
    fabric_mrepair_fuse_rbact2_i                             : in std_logic;
    fabric_data_from_system_i                                : in std_logic;
    fabric_data_from_bist_i                                  : in std_logic_vector(23 downto 0);
    fabric_otp_apb_enable_i                                  : in std_logic;
    fabric_mrepair_fuse_tm_i                                 : in std_logic;
    fabric_otp_security_rbact2_i                             : in std_logic;
    fabric_otp_security_rbact1_i                             : in std_logic;
    fabric_shift_en_i                                        : in std_logic_vector(23 downto 0);
    fabric_otp_cfg_loader_write_en_i                         : in std_logic;
    fabric_user_data_i                                       : in std_logic_vector(31 downto 0);
    fabric_mrepair_fuse_suppadd_i                            : in std_logic;
    fabric_mrepair_fuse_prog_i                               : in std_logic;
    fabric_otp_user_wordlock_i                               : in std_logic;
    fabric_ahb_direct_data_i                                 : in std_logic_vector(31 downto 0);
    fabric_otp_user_prog_i                                   : in std_logic;
    fabric_pd_active_i                                       : in std_logic_vector(23 downto 0);
    fabric_otp_user_suppadd_i                                : in std_logic;
    fabric_mrepair_fuse_pdn_i                                : in std_logic;
    fabric_otp_security_scanin_i                             : in std_logic_vector(4 downto 0);
    fabric_end_encoding_i                                    : in std_logic;
    fabric_jtag_tdo_usr2_i                                   : in std_logic;
    fabric_mrepair_fuse_wordlock_i                           : in std_logic;
    fabric_otp_user_prgwidth_i                               : in std_logic_vector(2 downto 0);
    fabric_otp_user_read_i                                   : in std_logic;
    fabric_mrepair_fuse_add_i                                : in std_logic_vector(6 downto 0);
    fabric_mrepair_fuse_bistmode_i                           : in std_logic;
    fabric_jtag_tdo_usr1_i                                   : in std_logic;
    fabric_otp_cfg_clk_fab_en_i                              : in std_logic;
    fabric_io_in_i                                           : in std_logic_vector(24 downto 0);
    fabric_sif_load_en_i                                     : in std_logic_vector(23 downto 0);
    fabric_mrepair_fuse_din_i                                : in std_logic_vector(38 downto 0);
    fabric_otp_apb_addr_i                                    : in std_logic_vector(31 downto 0);
    fabric_otp_apb_sel_i                                     : in std_logic;
    fabric_mrepair_fuse_rbact1_i                             : in std_logic;
    fabric_mrepair_fuse_configreg_i                          : in std_logic_vector(31 downto 0);
    fabric_otp_cfg_fabric_apb_en_i                           : in std_logic;
    fabric_data_shift_en_i                                   : in std_logic;
    fabric_lowskew_i21                                       : in std_logic;
    fabric_direct_data_i                                     : in std_logic_vector(31 downto 0);
    fabric_otp_user_pdn_i                                    : in std_logic;
    fabric_io_oe_i                                           : in std_logic_vector(24 downto 0);
    fabric_parusr_data_i                                     : in std_logic_vector(15 downto 0);
    fabric_otp_apb_write_i                                   : in std_logic;
    fabric_otp_security_testmode_i                           : in std_logic;
    fabric_system_data_to_mem_bist_i                         : in std_logic_vector(23 downto 0);
    fabric_tst_atpg_mrepair_i                                : in std_logic;
    fabric_mrepair_fuse_tstscanenable_i                      : in std_logic;
    fabric_otp_security_bistmode_i                           : in std_logic;
    fabric_lowskew_i22                                       : in std_logic;
    fabric_lowskew_i23                                       : in std_logic;
    fabric_lowskew_i20                                       : in std_logic;
    fabric_otp_user_configreg_i                              : in std_logic_vector(31 downto 0);
    fabric_otp_user_tst_scanin_i                             : in std_logic_vector(4 downto 0);
    fabric_sif_update_en_i                                   : in std_logic_vector(23 downto 0);
    fabric_mrepair_por_i                                     : in std_logic;
    fabric_mrepair_rst_n_i                                   : in std_logic;
    fabric_mrepair_initn_i                                   : in std_logic;
    fabric_spare_i                                           : in std_logic_vector(2 downto 0);

    fabric_mrepair_fuse_bbad_o                               : out std_logic;
    fabric_jtag_trst_n_o                                     : out std_logic;
    fabric_debug_direct_permission_write_o                   : out std_logic_vector(3 downto 0);
    fabric_otp_security_bist_end1_o                          : out std_logic;
    fabric_parusr_data_val_o                                 : out std_logic;
    fabric_debug_lock_reg_o                                  : out std_logic;
    fabric_debug_security_error_read_o                       : out std_logic;
    fabric_mrepair_fuse_tstscanout_o                         : out std_logic_vector(4 downto 0);
    fabric_otp_user_tst_scanout_o                            : out std_logic_vector(4 downto 0);
    fabric_sif_update_en_to_bist_o                           : out std_logic_vector(23 downto 0);
    fabric_otp_user_locked_o                                 : out std_logic;
    fabric_otp_security_bist_bad_o                           : out std_logic;
    fabric_debug_frame_permission_frame_o                    : out std_logic_vector(3 downto 0);
    fabric_otp_user_pwok_o                                   : out std_logic;
    fabric_otp_user_bend2_o                                  : out std_logic;
    fabric_mrepair_fuse_ded_o                                : out std_logic;
    fabric_debug_access_reg_data_ready_o                     : out std_logic;
    fabric_data_to_bist_o                                    : out std_logic_vector(23 downto 0);
    fabric_otp_user_startword_o                              : out std_logic_vector(15 downto 0);
    fabric_ahb_direct_data_o                                 : out std_logic_vector(31 downto 0);
    fabric_parusr_data_o                                     : out std_logic_vector(15 downto 0);
    fabric_debug_otp_reload_err_o                            : out std_logic;
    fabric_cfg_fabric_user_unmask_o                          : out std_logic;
    fabric_decoder_init_ready_o                              : out std_logic;
    fabric_global_chip_status_o                              : out std_logic_vector(2 downto 0);
    fabric_debug_security_boot_done_o                        : out std_logic;
    fabric_otp_user_calibrated_o                             : out std_logic;
    fabric_fuse_status_o                                     : out std_logic_vector(2 downto 0);
    fabric_otp_apb_rdata_o                                   : out std_logic_vector(31 downto 0);
    fabric_jtag_tms_o                                        : out std_logic;
    fabric_debug_bsec_core_status_o                          : out std_logic_vector(31 downto 0);
    fabric_mrepair_fuse_bist1fail_o                          : out std_logic_vector(7 downto 0);
    fabric_flag_ready_o                                      : out std_logic;
    fabric_mrepair_fuse_dout_o                               : out std_logic_vector(40 downto 0);
    fabric_debug_rst_soft_o                                  : out std_logic;
    fabric_otp_user_ack_o                                    : out std_logic;
    fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o  : out std_logic;
    fabric_shift_en_to_bist_o                                : out std_logic_vector(23 downto 0);
    fabric_sif_reg_en_to_bist_o                              : out std_logic_vector(119 downto 0);
    fabric_debug_otp_manager_read_otp_o                      : out std_logic;
    fabric_otp_user_sec_o                                    : out std_logic;
    fabric_otp_user_wlromout_o                               : out std_logic_vector(9 downto 0);
    fabric_mrepair_fuse_bend1_o                              : out std_logic;
    fabric_mrepair_fuse_flagstate_o                          : out std_logic_vector(3 downto 0);
    fabric_system_data_from_mem_bist_o                       : out std_logic_vector(23 downto 0);
    fabric_direct_data_o                                     : out std_logic_vector(31 downto 0);
    fabric_otp_user_bbad_o                                   : out std_logic;
    fabric_user_read_cycle_o                                 : out std_logic;
    fabric_chip_status_o                                     : out std_logic_vector(71 downto 0);
    fabric_mrepair_fuse_disturbed_o                          : out std_logic;
    fabric_debug_otpboot_state_o                             : out std_logic_vector(2 downto 0);
    fabric_pd_ready_o                                        : out std_logic_vector(23 downto 0);
    fabric_debug_key_correct_o                               : out std_logic;
    fabric_otp_apb_ready_o                                   : out std_logic;
    fabric_otp_user_progfail_o                               : out std_logic;
    fabric_mrepair_fuse_sec_o                                : out std_logic;
    fabric_mrepair_fuse_bend2_o                              : out std_logic;
    fabric_debug_lifecycle_o                                 : out std_logic_vector(3 downto 0);
    fabric_mrepair_fuse_ack_o                                : out std_logic;
    fabric_debug_cpt_retry_o                                 : out std_logic_vector(3 downto 0);
    fabric_otp_security_ack_o                                : out std_logic;
    fabric_debug_otpmgmt_state_o                             : out std_logic_vector(2 downto 0);
    fabric_mrepair_fuse_progfail_o                           : out std_logic;
    fabric_otp_user_bist2fail_o                              : out std_logic_vector(6 downto 0);
    fabric_user_data_o                                       : out std_logic_vector(31 downto 0);
    fabric_jtag_tdi_o                                        : out std_logic;
    fabric_lowskew_o3                                        : out std_logic;
    fabric_lowskew_o5                                        : out std_logic;
    fabric_lowskew_o4                                        : out std_logic;
    fabric_debug_error_o                                     : out std_logic;
    fabric_jtag_usr2_o                                       : out std_logic;
    fabric_mrepair_fuse_wlromout_o                           : out std_logic_vector(9 downto 0);
    fabric_debug_otpapb_state_o                              : out std_logic_vector(2 downto 0);
    fabric_otp_user_bist1fail_o                              : out std_logic_vector(7 downto 0);
    fabric_otp_security_bist_fail2_o                         : out std_logic_vector(6 downto 0);
    fabric_otp_user_disturbed_o                              : out std_logic;
    fabric_flag_trigger_o                                    : out std_logic;
    fabric_otp_security_bist_end2_o                          : out std_logic;
    fabric_otp_security_bist_fail1_o                         : out std_logic_vector(7 downto 0);
    fabric_mrepair_fuse_locked_o                             : out std_logic;
    fabric_otp_user_flagstate_o                              : out std_logic_vector(3 downto 0);
    fabric_otp_security_scanout_o                            : out std_logic_vector(4 downto 0);
    fabric_user_write_cycle_o                                : out std_logic;
    fabric_debug_fsm_state_o                                 : out std_logic_vector(2 downto 0);
    fabric_otp_user_ded_o                                    : out std_logic;
    fabric_debug_otp_manager_read_done_o                     : out std_logic;
    fabric_debug_frame_use_encryption_o                      : out std_logic;
    fabric_data_to_system_o                                  : out std_logic;
    fabric_jtag_usr1_o                                       : out std_logic;
    fabric_otp_user_bend1_o                                  : out std_logic;
    fabric_debug_otpboot_curr_addr_o                         : out std_logic_vector(7 downto 0);
    fabric_mrepair_fuse_ready_o                              : out std_logic;
    fabric_mrepair_fuse_calibrated_o                         : out std_logic;
    fabric_sif_load_en_to_bist_o                             : out std_logic_vector(23 downto 0);
    fabric_io_out_o                                          : out std_logic_vector(24 downto 0);
    fabric_mrepair_fuse_startword_o                          : out std_logic_vector(15 downto 0);
    fabric_system_dataready_o                                : out std_logic;
    fabric_mrepair_fuse_pwok_o                               : out std_logic;
    fabric_lowskew_o6                                        : out std_logic;
    fabric_cfg_fabric_user_flag_o                            : out std_logic;
    fabric_otp_user_dout_o                                   : out std_logic_vector(40 downto 0);
    fabric_mrepair_fuse_bist2fail_o                          : out std_logic_vector(6 downto 0);
    fabric_status_cold_start_o                               : out std_logic;
    fabric_flag_error_o                                      : out std_logic;
    fabric_debug_direct_permission_read_o                    : out std_logic_vector(3 downto 0)
);
end NX_SERVICE_U_WRAP;

architecture NX_ARCH of NX_SERVICE_U_WRAP is
begin

    inst_NX_SERVICE_U : NX_SERVICE_U
    generic map (
         bsm_config                                                => bsm_config
       , ahb_config                                                => ahb_config
    )
    port map (
         fabric_otp_user_tst_scanenable_i                         => fabric_otp_user_tst_scanenable_i
       , fabric_otp_cfg_loader_read_en_i                          => fabric_otp_cfg_loader_read_en_i
       , fabric_otp_security_force_pdn1_i                         => fabric_otp_security_force_pdn1_i
       , fabric_otp_security_scanenable_i                         => fabric_otp_security_scanenable_i
       , fabric_otp_user_din_i1                                   => fabric_otp_user_din_i(0)
       , fabric_otp_user_din_i2                                   => fabric_otp_user_din_i(1)
       , fabric_otp_user_din_i3                                   => fabric_otp_user_din_i(2)
       , fabric_otp_user_din_i4                                   => fabric_otp_user_din_i(3)
       , fabric_otp_user_din_i5                                   => fabric_otp_user_din_i(4)
       , fabric_otp_user_din_i6                                   => fabric_otp_user_din_i(5)
       , fabric_otp_user_din_i7                                   => fabric_otp_user_din_i(6)
       , fabric_otp_user_din_i8                                   => fabric_otp_user_din_i(7)
       , fabric_otp_user_din_i9                                   => fabric_otp_user_din_i(8)
       , fabric_otp_user_din_i10                                  => fabric_otp_user_din_i(9)
       , fabric_otp_user_din_i11                                  => fabric_otp_user_din_i(10)
       , fabric_otp_user_din_i12                                  => fabric_otp_user_din_i(11)
       , fabric_otp_user_din_i13                                  => fabric_otp_user_din_i(12)
       , fabric_otp_user_din_i14                                  => fabric_otp_user_din_i(13)
       , fabric_otp_user_din_i15                                  => fabric_otp_user_din_i(14)
       , fabric_otp_user_din_i16                                  => fabric_otp_user_din_i(15)
       , fabric_otp_user_din_i17                                  => fabric_otp_user_din_i(16)
       , fabric_otp_user_din_i18                                  => fabric_otp_user_din_i(17)
       , fabric_otp_user_din_i19                                  => fabric_otp_user_din_i(18)
       , fabric_otp_user_din_i20                                  => fabric_otp_user_din_i(19)
       , fabric_otp_user_din_i21                                  => fabric_otp_user_din_i(20)
       , fabric_otp_user_din_i22                                  => fabric_otp_user_din_i(21)
       , fabric_otp_user_din_i23                                  => fabric_otp_user_din_i(22)
       , fabric_otp_user_din_i24                                  => fabric_otp_user_din_i(23)
       , fabric_otp_user_din_i25                                  => fabric_otp_user_din_i(24)
       , fabric_otp_user_din_i26                                  => fabric_otp_user_din_i(25)
       , fabric_otp_user_din_i27                                  => fabric_otp_user_din_i(26)
       , fabric_otp_user_din_i28                                  => fabric_otp_user_din_i(27)
       , fabric_otp_user_din_i29                                  => fabric_otp_user_din_i(28)
       , fabric_otp_user_din_i30                                  => fabric_otp_user_din_i(29)
       , fabric_otp_user_din_i31                                  => fabric_otp_user_din_i(30)
       , fabric_otp_user_din_i32                                  => fabric_otp_user_din_i(31)
       , fabric_otp_user_din_i33                                  => fabric_otp_user_din_i(32)
       , fabric_otp_user_din_i34                                  => fabric_otp_user_din_i(33)
       , fabric_otp_user_din_i35                                  => fabric_otp_user_din_i(34)
       , fabric_otp_user_din_i36                                  => fabric_otp_user_din_i(35)
       , fabric_otp_user_din_i37                                  => fabric_otp_user_din_i(36)
       , fabric_otp_user_din_i38                                  => fabric_otp_user_din_i(37)
       , fabric_otp_user_din_i39                                  => fabric_otp_user_din_i(38)
       , fabric_mrepair_fuse_prgwidth_i1                          => fabric_mrepair_fuse_prgwidth_i(0)
       , fabric_mrepair_fuse_prgwidth_i2                          => fabric_mrepair_fuse_prgwidth_i(1)
       , fabric_mrepair_fuse_prgwidth_i3                          => fabric_mrepair_fuse_prgwidth_i(2)
       , fabric_otp_apb_wdata_i1                                  => fabric_otp_apb_wdata_i(0)
       , fabric_otp_apb_wdata_i2                                  => fabric_otp_apb_wdata_i(1)
       , fabric_otp_apb_wdata_i3                                  => fabric_otp_apb_wdata_i(2)
       , fabric_otp_apb_wdata_i4                                  => fabric_otp_apb_wdata_i(3)
       , fabric_otp_apb_wdata_i5                                  => fabric_otp_apb_wdata_i(4)
       , fabric_otp_apb_wdata_i6                                  => fabric_otp_apb_wdata_i(5)
       , fabric_otp_apb_wdata_i7                                  => fabric_otp_apb_wdata_i(6)
       , fabric_otp_apb_wdata_i8                                  => fabric_otp_apb_wdata_i(7)
       , fabric_otp_apb_wdata_i9                                  => fabric_otp_apb_wdata_i(8)
       , fabric_otp_apb_wdata_i10                                 => fabric_otp_apb_wdata_i(9)
       , fabric_otp_apb_wdata_i11                                 => fabric_otp_apb_wdata_i(10)
       , fabric_otp_apb_wdata_i12                                 => fabric_otp_apb_wdata_i(11)
       , fabric_otp_apb_wdata_i13                                 => fabric_otp_apb_wdata_i(12)
       , fabric_otp_apb_wdata_i14                                 => fabric_otp_apb_wdata_i(13)
       , fabric_otp_apb_wdata_i15                                 => fabric_otp_apb_wdata_i(14)
       , fabric_otp_apb_wdata_i16                                 => fabric_otp_apb_wdata_i(15)
       , fabric_otp_apb_wdata_i17                                 => fabric_otp_apb_wdata_i(16)
       , fabric_otp_apb_wdata_i18                                 => fabric_otp_apb_wdata_i(17)
       , fabric_otp_apb_wdata_i19                                 => fabric_otp_apb_wdata_i(18)
       , fabric_otp_apb_wdata_i20                                 => fabric_otp_apb_wdata_i(19)
       , fabric_otp_apb_wdata_i21                                 => fabric_otp_apb_wdata_i(20)
       , fabric_otp_apb_wdata_i22                                 => fabric_otp_apb_wdata_i(21)
       , fabric_otp_apb_wdata_i23                                 => fabric_otp_apb_wdata_i(22)
       , fabric_otp_apb_wdata_i24                                 => fabric_otp_apb_wdata_i(23)
       , fabric_otp_apb_wdata_i25                                 => fabric_otp_apb_wdata_i(24)
       , fabric_otp_apb_wdata_i26                                 => fabric_otp_apb_wdata_i(25)
       , fabric_otp_apb_wdata_i27                                 => fabric_otp_apb_wdata_i(26)
       , fabric_otp_apb_wdata_i28                                 => fabric_otp_apb_wdata_i(27)
       , fabric_otp_apb_wdata_i29                                 => fabric_otp_apb_wdata_i(28)
       , fabric_otp_apb_wdata_i30                                 => fabric_otp_apb_wdata_i(29)
       , fabric_otp_apb_wdata_i31                                 => fabric_otp_apb_wdata_i(30)
       , fabric_otp_apb_wdata_i32                                 => fabric_otp_apb_wdata_i(31)
       , fabric_otp_cfg_clk_otpm_disable_i                        => fabric_otp_cfg_clk_otpm_disable_i
       , fabric_otp_user_disturbcheck_i                           => fabric_otp_user_disturbcheck_i
       , fabric_mrepair_fuse_read_i                               => fabric_mrepair_fuse_read_i
       , fabric_otp_user_rbact2_i                                 => fabric_otp_user_rbact2_i
       , fabric_mrepair_fuse_eccbypass_i                          => fabric_mrepair_fuse_eccbypass_i
       , fabric_otp_user_bistmode_i                               => fabric_otp_user_bistmode_i
       , fabric_otp_user_add_i1                                   => fabric_otp_user_add_i(0)
       , fabric_otp_user_add_i2                                   => fabric_otp_user_add_i(1)
       , fabric_otp_user_add_i3                                   => fabric_otp_user_add_i(2)
       , fabric_otp_user_add_i4                                   => fabric_otp_user_add_i(3)
       , fabric_otp_user_add_i5                                   => fabric_otp_user_add_i(4)
       , fabric_otp_user_add_i6                                   => fabric_otp_user_add_i(5)
       , fabric_otp_user_add_i7                                   => fabric_otp_user_add_i(6)
       , fabric_otp_user_tm_i                                     => fabric_otp_user_tm_i
       , fabric_otp_rstn_i                                        => fabric_otp_rstn_i
       , fabric_mrepair_fuse_disturbchecked_i                     => fabric_mrepair_fuse_disturbchecked_i
       , fabric_otp_user_rbact1_i                                 => fabric_otp_user_rbact1_i
       , fabric_mrepair_fuse_tst_scanin_i1                        => fabric_mrepair_fuse_tst_scanin_i(0)
       , fabric_mrepair_fuse_tst_scanin_i2                        => fabric_mrepair_fuse_tst_scanin_i(1)
       , fabric_mrepair_fuse_tst_scanin_i3                        => fabric_mrepair_fuse_tst_scanin_i(2)
       , fabric_mrepair_fuse_tst_scanin_i4                        => fabric_mrepair_fuse_tst_scanin_i(3)
       , fabric_mrepair_fuse_tst_scanin_i5                        => fabric_mrepair_fuse_tst_scanin_i(4)
       , fabric_parusr_type_i1                                    => fabric_parusr_type_i(0)
       , fabric_parusr_type_i2                                    => fabric_parusr_type_i(1)
       , fabric_mrepair_fuse_redbypass_i                          => fabric_mrepair_fuse_redbypass_i
       , fabric_otp_user_eccbypass_i                              => fabric_otp_user_eccbypass_i
       , fabric_otp_user_redbypass_i                              => fabric_otp_user_redbypass_i
       , fabric_mrepair_mode_i1                                   => fabric_mrepair_mode_i(0)
       , fabric_mrepair_mode_i2                                   => fabric_mrepair_mode_i(1)
       , fabric_mrepair_mode_i3                                   => fabric_mrepair_mode_i(2)
       , fabric_mrepair_mode_i4                                   => fabric_mrepair_mode_i(3)
       , fabric_parusr_cs_i                                       => fabric_parusr_cs_i
       , fabric_sif_reg_en_i1                                     => fabric_sif_reg_en_i(0)
       , fabric_sif_reg_en_i2                                     => fabric_sif_reg_en_i(1)
       , fabric_sif_reg_en_i3                                     => fabric_sif_reg_en_i(2)
       , fabric_sif_reg_en_i4                                     => fabric_sif_reg_en_i(3)
       , fabric_sif_reg_en_i5                                     => fabric_sif_reg_en_i(4)
       , fabric_sif_reg_en_i6                                     => fabric_sif_reg_en_i(5)
       , fabric_sif_reg_en_i7                                     => fabric_sif_reg_en_i(6)
       , fabric_sif_reg_en_i8                                     => fabric_sif_reg_en_i(7)
       , fabric_sif_reg_en_i9                                     => fabric_sif_reg_en_i(8)
       , fabric_sif_reg_en_i10                                    => fabric_sif_reg_en_i(9)
       , fabric_sif_reg_en_i11                                    => fabric_sif_reg_en_i(10)
       , fabric_sif_reg_en_i12                                    => fabric_sif_reg_en_i(11)
       , fabric_sif_reg_en_i13                                    => fabric_sif_reg_en_i(12)
       , fabric_sif_reg_en_i14                                    => fabric_sif_reg_en_i(13)
       , fabric_sif_reg_en_i15                                    => fabric_sif_reg_en_i(14)
       , fabric_sif_reg_en_i16                                    => fabric_sif_reg_en_i(15)
       , fabric_sif_reg_en_i17                                    => fabric_sif_reg_en_i(16)
       , fabric_sif_reg_en_i18                                    => fabric_sif_reg_en_i(17)
       , fabric_sif_reg_en_i19                                    => fabric_sif_reg_en_i(18)
       , fabric_sif_reg_en_i20                                    => fabric_sif_reg_en_i(19)
       , fabric_sif_reg_en_i21                                    => fabric_sif_reg_en_i(20)
       , fabric_sif_reg_en_i22                                    => fabric_sif_reg_en_i(21)
       , fabric_sif_reg_en_i23                                    => fabric_sif_reg_en_i(22)
       , fabric_sif_reg_en_i24                                    => fabric_sif_reg_en_i(23)
       , fabric_sif_reg_en_i25                                    => fabric_sif_reg_en_i(24)
       , fabric_sif_reg_en_i26                                    => fabric_sif_reg_en_i(25)
       , fabric_sif_reg_en_i27                                    => fabric_sif_reg_en_i(26)
       , fabric_sif_reg_en_i28                                    => fabric_sif_reg_en_i(27)
       , fabric_sif_reg_en_i29                                    => fabric_sif_reg_en_i(28)
       , fabric_sif_reg_en_i30                                    => fabric_sif_reg_en_i(29)
       , fabric_sif_reg_en_i31                                    => fabric_sif_reg_en_i(30)
       , fabric_sif_reg_en_i32                                    => fabric_sif_reg_en_i(31)
       , fabric_sif_reg_en_i33                                    => fabric_sif_reg_en_i(32)
       , fabric_sif_reg_en_i34                                    => fabric_sif_reg_en_i(33)
       , fabric_sif_reg_en_i35                                    => fabric_sif_reg_en_i(34)
       , fabric_sif_reg_en_i36                                    => fabric_sif_reg_en_i(35)
       , fabric_sif_reg_en_i37                                    => fabric_sif_reg_en_i(36)
       , fabric_sif_reg_en_i38                                    => fabric_sif_reg_en_i(37)
       , fabric_sif_reg_en_i39                                    => fabric_sif_reg_en_i(38)
       , fabric_sif_reg_en_i40                                    => fabric_sif_reg_en_i(39)
       , fabric_sif_reg_en_i41                                    => fabric_sif_reg_en_i(40)
       , fabric_sif_reg_en_i42                                    => fabric_sif_reg_en_i(41)
       , fabric_sif_reg_en_i43                                    => fabric_sif_reg_en_i(42)
       , fabric_sif_reg_en_i44                                    => fabric_sif_reg_en_i(43)
       , fabric_sif_reg_en_i45                                    => fabric_sif_reg_en_i(44)
       , fabric_sif_reg_en_i46                                    => fabric_sif_reg_en_i(45)
       , fabric_sif_reg_en_i47                                    => fabric_sif_reg_en_i(46)
       , fabric_sif_reg_en_i48                                    => fabric_sif_reg_en_i(47)
       , fabric_sif_reg_en_i49                                    => fabric_sif_reg_en_i(48)
       , fabric_sif_reg_en_i50                                    => fabric_sif_reg_en_i(49)
       , fabric_sif_reg_en_i51                                    => fabric_sif_reg_en_i(50)
       , fabric_sif_reg_en_i52                                    => fabric_sif_reg_en_i(51)
       , fabric_sif_reg_en_i53                                    => fabric_sif_reg_en_i(52)
       , fabric_sif_reg_en_i54                                    => fabric_sif_reg_en_i(53)
       , fabric_sif_reg_en_i55                                    => fabric_sif_reg_en_i(54)
       , fabric_sif_reg_en_i56                                    => fabric_sif_reg_en_i(55)
       , fabric_sif_reg_en_i57                                    => fabric_sif_reg_en_i(56)
       , fabric_sif_reg_en_i58                                    => fabric_sif_reg_en_i(57)
       , fabric_sif_reg_en_i59                                    => fabric_sif_reg_en_i(58)
       , fabric_sif_reg_en_i60                                    => fabric_sif_reg_en_i(59)
       , fabric_sif_reg_en_i61                                    => fabric_sif_reg_en_i(60)
       , fabric_sif_reg_en_i62                                    => fabric_sif_reg_en_i(61)
       , fabric_sif_reg_en_i63                                    => fabric_sif_reg_en_i(62)
       , fabric_sif_reg_en_i64                                    => fabric_sif_reg_en_i(63)
       , fabric_sif_reg_en_i65                                    => fabric_sif_reg_en_i(64)
       , fabric_sif_reg_en_i66                                    => fabric_sif_reg_en_i(65)
       , fabric_sif_reg_en_i67                                    => fabric_sif_reg_en_i(66)
       , fabric_sif_reg_en_i68                                    => fabric_sif_reg_en_i(67)
       , fabric_sif_reg_en_i69                                    => fabric_sif_reg_en_i(68)
       , fabric_sif_reg_en_i70                                    => fabric_sif_reg_en_i(69)
       , fabric_sif_reg_en_i71                                    => fabric_sif_reg_en_i(70)
       , fabric_sif_reg_en_i72                                    => fabric_sif_reg_en_i(71)
       , fabric_sif_reg_en_i73                                    => fabric_sif_reg_en_i(72)
       , fabric_sif_reg_en_i74                                    => fabric_sif_reg_en_i(73)
       , fabric_sif_reg_en_i75                                    => fabric_sif_reg_en_i(74)
       , fabric_sif_reg_en_i76                                    => fabric_sif_reg_en_i(75)
       , fabric_sif_reg_en_i77                                    => fabric_sif_reg_en_i(76)
       , fabric_sif_reg_en_i78                                    => fabric_sif_reg_en_i(77)
       , fabric_sif_reg_en_i79                                    => fabric_sif_reg_en_i(78)
       , fabric_sif_reg_en_i80                                    => fabric_sif_reg_en_i(79)
       , fabric_sif_reg_en_i81                                    => fabric_sif_reg_en_i(80)
       , fabric_sif_reg_en_i82                                    => fabric_sif_reg_en_i(81)
       , fabric_sif_reg_en_i83                                    => fabric_sif_reg_en_i(82)
       , fabric_sif_reg_en_i84                                    => fabric_sif_reg_en_i(83)
       , fabric_sif_reg_en_i85                                    => fabric_sif_reg_en_i(84)
       , fabric_sif_reg_en_i86                                    => fabric_sif_reg_en_i(85)
       , fabric_sif_reg_en_i87                                    => fabric_sif_reg_en_i(86)
       , fabric_sif_reg_en_i88                                    => fabric_sif_reg_en_i(87)
       , fabric_sif_reg_en_i89                                    => fabric_sif_reg_en_i(88)
       , fabric_sif_reg_en_i90                                    => fabric_sif_reg_en_i(89)
       , fabric_sif_reg_en_i91                                    => fabric_sif_reg_en_i(90)
       , fabric_sif_reg_en_i92                                    => fabric_sif_reg_en_i(91)
       , fabric_sif_reg_en_i93                                    => fabric_sif_reg_en_i(92)
       , fabric_sif_reg_en_i94                                    => fabric_sif_reg_en_i(93)
       , fabric_sif_reg_en_i95                                    => fabric_sif_reg_en_i(94)
       , fabric_sif_reg_en_i96                                    => fabric_sif_reg_en_i(95)
       , fabric_sif_reg_en_i97                                    => fabric_sif_reg_en_i(96)
       , fabric_sif_reg_en_i98                                    => fabric_sif_reg_en_i(97)
       , fabric_sif_reg_en_i99                                    => fabric_sif_reg_en_i(98)
       , fabric_sif_reg_en_i100                                   => fabric_sif_reg_en_i(99)
       , fabric_sif_reg_en_i101                                   => fabric_sif_reg_en_i(100)
       , fabric_sif_reg_en_i102                                   => fabric_sif_reg_en_i(101)
       , fabric_sif_reg_en_i103                                   => fabric_sif_reg_en_i(102)
       , fabric_sif_reg_en_i104                                   => fabric_sif_reg_en_i(103)
       , fabric_sif_reg_en_i105                                   => fabric_sif_reg_en_i(104)
       , fabric_sif_reg_en_i106                                   => fabric_sif_reg_en_i(105)
       , fabric_sif_reg_en_i107                                   => fabric_sif_reg_en_i(106)
       , fabric_sif_reg_en_i108                                   => fabric_sif_reg_en_i(107)
       , fabric_sif_reg_en_i109                                   => fabric_sif_reg_en_i(108)
       , fabric_sif_reg_en_i110                                   => fabric_sif_reg_en_i(109)
       , fabric_sif_reg_en_i111                                   => fabric_sif_reg_en_i(110)
       , fabric_sif_reg_en_i112                                   => fabric_sif_reg_en_i(111)
       , fabric_sif_reg_en_i113                                   => fabric_sif_reg_en_i(112)
       , fabric_sif_reg_en_i114                                   => fabric_sif_reg_en_i(113)
       , fabric_sif_reg_en_i115                                   => fabric_sif_reg_en_i(114)
       , fabric_sif_reg_en_i116                                   => fabric_sif_reg_en_i(115)
       , fabric_sif_reg_en_i117                                   => fabric_sif_reg_en_i(116)
       , fabric_sif_reg_en_i118                                   => fabric_sif_reg_en_i(117)
       , fabric_sif_reg_en_i119                                   => fabric_sif_reg_en_i(118)
       , fabric_sif_reg_en_i120                                   => fabric_sif_reg_en_i(119)
       , fabric_mrepair_fuse_rbact2_i                             => fabric_mrepair_fuse_rbact2_i
       , fabric_data_from_system_i                                => fabric_data_from_system_i
       , fabric_data_from_bist_i1                                 => fabric_data_from_bist_i(0)
       , fabric_data_from_bist_i2                                 => fabric_data_from_bist_i(1)
       , fabric_data_from_bist_i3                                 => fabric_data_from_bist_i(2)
       , fabric_data_from_bist_i4                                 => fabric_data_from_bist_i(3)
       , fabric_data_from_bist_i5                                 => fabric_data_from_bist_i(4)
       , fabric_data_from_bist_i6                                 => fabric_data_from_bist_i(5)
       , fabric_data_from_bist_i7                                 => fabric_data_from_bist_i(6)
       , fabric_data_from_bist_i8                                 => fabric_data_from_bist_i(7)
       , fabric_data_from_bist_i9                                 => fabric_data_from_bist_i(8)
       , fabric_data_from_bist_i10                                => fabric_data_from_bist_i(9)
       , fabric_data_from_bist_i11                                => fabric_data_from_bist_i(10)
       , fabric_data_from_bist_i12                                => fabric_data_from_bist_i(11)
       , fabric_data_from_bist_i13                                => fabric_data_from_bist_i(12)
       , fabric_data_from_bist_i14                                => fabric_data_from_bist_i(13)
       , fabric_data_from_bist_i15                                => fabric_data_from_bist_i(14)
       , fabric_data_from_bist_i16                                => fabric_data_from_bist_i(15)
       , fabric_data_from_bist_i17                                => fabric_data_from_bist_i(16)
       , fabric_data_from_bist_i18                                => fabric_data_from_bist_i(17)
       , fabric_data_from_bist_i19                                => fabric_data_from_bist_i(18)
       , fabric_data_from_bist_i20                                => fabric_data_from_bist_i(19)
       , fabric_data_from_bist_i21                                => fabric_data_from_bist_i(20)
       , fabric_data_from_bist_i22                                => fabric_data_from_bist_i(21)
       , fabric_data_from_bist_i23                                => fabric_data_from_bist_i(22)
       , fabric_data_from_bist_i24                                => fabric_data_from_bist_i(23)
       , fabric_otp_apb_enable_i                                  => fabric_otp_apb_enable_i
       , fabric_mrepair_fuse_tm_i                                 => fabric_mrepair_fuse_tm_i
       , fabric_otp_security_rbact2_i                             => fabric_otp_security_rbact2_i
       , fabric_otp_security_rbact1_i                             => fabric_otp_security_rbact1_i
       , fabric_shift_en_i1                                       => fabric_shift_en_i(0)
       , fabric_shift_en_i2                                       => fabric_shift_en_i(1)
       , fabric_shift_en_i3                                       => fabric_shift_en_i(2)
       , fabric_shift_en_i4                                       => fabric_shift_en_i(3)
       , fabric_shift_en_i5                                       => fabric_shift_en_i(4)
       , fabric_shift_en_i6                                       => fabric_shift_en_i(5)
       , fabric_shift_en_i7                                       => fabric_shift_en_i(6)
       , fabric_shift_en_i8                                       => fabric_shift_en_i(7)
       , fabric_shift_en_i9                                       => fabric_shift_en_i(8)
       , fabric_shift_en_i10                                      => fabric_shift_en_i(9)
       , fabric_shift_en_i11                                      => fabric_shift_en_i(10)
       , fabric_shift_en_i12                                      => fabric_shift_en_i(11)
       , fabric_shift_en_i13                                      => fabric_shift_en_i(12)
       , fabric_shift_en_i14                                      => fabric_shift_en_i(13)
       , fabric_shift_en_i15                                      => fabric_shift_en_i(14)
       , fabric_shift_en_i16                                      => fabric_shift_en_i(15)
       , fabric_shift_en_i17                                      => fabric_shift_en_i(16)
       , fabric_shift_en_i18                                      => fabric_shift_en_i(17)
       , fabric_shift_en_i19                                      => fabric_shift_en_i(18)
       , fabric_shift_en_i20                                      => fabric_shift_en_i(19)
       , fabric_shift_en_i21                                      => fabric_shift_en_i(20)
       , fabric_shift_en_i22                                      => fabric_shift_en_i(21)
       , fabric_shift_en_i23                                      => fabric_shift_en_i(22)
       , fabric_shift_en_i24                                      => fabric_shift_en_i(23)
       , fabric_otp_cfg_loader_write_en_i                         => fabric_otp_cfg_loader_write_en_i
       , fabric_user_data_i1                                      => fabric_user_data_i(0)
       , fabric_user_data_i2                                      => fabric_user_data_i(1)
       , fabric_user_data_i3                                      => fabric_user_data_i(2)
       , fabric_user_data_i4                                      => fabric_user_data_i(3)
       , fabric_user_data_i5                                      => fabric_user_data_i(4)
       , fabric_user_data_i6                                      => fabric_user_data_i(5)
       , fabric_user_data_i7                                      => fabric_user_data_i(6)
       , fabric_user_data_i8                                      => fabric_user_data_i(7)
       , fabric_user_data_i9                                      => fabric_user_data_i(8)
       , fabric_user_data_i10                                     => fabric_user_data_i(9)
       , fabric_user_data_i11                                     => fabric_user_data_i(10)
       , fabric_user_data_i12                                     => fabric_user_data_i(11)
       , fabric_user_data_i13                                     => fabric_user_data_i(12)
       , fabric_user_data_i14                                     => fabric_user_data_i(13)
       , fabric_user_data_i15                                     => fabric_user_data_i(14)
       , fabric_user_data_i16                                     => fabric_user_data_i(15)
       , fabric_user_data_i17                                     => fabric_user_data_i(16)
       , fabric_user_data_i18                                     => fabric_user_data_i(17)
       , fabric_user_data_i19                                     => fabric_user_data_i(18)
       , fabric_user_data_i20                                     => fabric_user_data_i(19)
       , fabric_user_data_i21                                     => fabric_user_data_i(20)
       , fabric_user_data_i22                                     => fabric_user_data_i(21)
       , fabric_user_data_i23                                     => fabric_user_data_i(22)
       , fabric_user_data_i24                                     => fabric_user_data_i(23)
       , fabric_user_data_i25                                     => fabric_user_data_i(24)
       , fabric_user_data_i26                                     => fabric_user_data_i(25)
       , fabric_user_data_i27                                     => fabric_user_data_i(26)
       , fabric_user_data_i28                                     => fabric_user_data_i(27)
       , fabric_user_data_i29                                     => fabric_user_data_i(28)
       , fabric_user_data_i30                                     => fabric_user_data_i(29)
       , fabric_user_data_i31                                     => fabric_user_data_i(30)
       , fabric_user_data_i32                                     => fabric_user_data_i(31)
       , fabric_mrepair_fuse_suppadd_i                            => fabric_mrepair_fuse_suppadd_i
       , fabric_mrepair_fuse_prog_i                               => fabric_mrepair_fuse_prog_i
       , fabric_otp_user_wordlock_i                               => fabric_otp_user_wordlock_i
       , fabric_ahb_direct_data_i1                                => fabric_ahb_direct_data_i(0)
       , fabric_ahb_direct_data_i2                                => fabric_ahb_direct_data_i(1)
       , fabric_ahb_direct_data_i3                                => fabric_ahb_direct_data_i(2)
       , fabric_ahb_direct_data_i4                                => fabric_ahb_direct_data_i(3)
       , fabric_ahb_direct_data_i5                                => fabric_ahb_direct_data_i(4)
       , fabric_ahb_direct_data_i6                                => fabric_ahb_direct_data_i(5)
       , fabric_ahb_direct_data_i7                                => fabric_ahb_direct_data_i(6)
       , fabric_ahb_direct_data_i8                                => fabric_ahb_direct_data_i(7)
       , fabric_ahb_direct_data_i9                                => fabric_ahb_direct_data_i(8)
       , fabric_ahb_direct_data_i10                               => fabric_ahb_direct_data_i(9)
       , fabric_ahb_direct_data_i11                               => fabric_ahb_direct_data_i(10)
       , fabric_ahb_direct_data_i12                               => fabric_ahb_direct_data_i(11)
       , fabric_ahb_direct_data_i13                               => fabric_ahb_direct_data_i(12)
       , fabric_ahb_direct_data_i14                               => fabric_ahb_direct_data_i(13)
       , fabric_ahb_direct_data_i15                               => fabric_ahb_direct_data_i(14)
       , fabric_ahb_direct_data_i16                               => fabric_ahb_direct_data_i(15)
       , fabric_ahb_direct_data_i17                               => fabric_ahb_direct_data_i(16)
       , fabric_ahb_direct_data_i18                               => fabric_ahb_direct_data_i(17)
       , fabric_ahb_direct_data_i19                               => fabric_ahb_direct_data_i(18)
       , fabric_ahb_direct_data_i20                               => fabric_ahb_direct_data_i(19)
       , fabric_ahb_direct_data_i21                               => fabric_ahb_direct_data_i(20)
       , fabric_ahb_direct_data_i22                               => fabric_ahb_direct_data_i(21)
       , fabric_ahb_direct_data_i23                               => fabric_ahb_direct_data_i(22)
       , fabric_ahb_direct_data_i24                               => fabric_ahb_direct_data_i(23)
       , fabric_ahb_direct_data_i25                               => fabric_ahb_direct_data_i(24)
       , fabric_ahb_direct_data_i26                               => fabric_ahb_direct_data_i(25)
       , fabric_ahb_direct_data_i27                               => fabric_ahb_direct_data_i(26)
       , fabric_ahb_direct_data_i28                               => fabric_ahb_direct_data_i(27)
       , fabric_ahb_direct_data_i29                               => fabric_ahb_direct_data_i(28)
       , fabric_ahb_direct_data_i30                               => fabric_ahb_direct_data_i(29)
       , fabric_ahb_direct_data_i31                               => fabric_ahb_direct_data_i(30)
       , fabric_ahb_direct_data_i32                               => fabric_ahb_direct_data_i(31)
       , fabric_otp_user_prog_i                                   => fabric_otp_user_prog_i
       , fabric_pd_active_i1                                      => fabric_pd_active_i(0)
       , fabric_pd_active_i2                                      => fabric_pd_active_i(1)
       , fabric_pd_active_i3                                      => fabric_pd_active_i(2)
       , fabric_pd_active_i4                                      => fabric_pd_active_i(3)
       , fabric_pd_active_i5                                      => fabric_pd_active_i(4)
       , fabric_pd_active_i6                                      => fabric_pd_active_i(5)
       , fabric_pd_active_i7                                      => fabric_pd_active_i(6)
       , fabric_pd_active_i8                                      => fabric_pd_active_i(7)
       , fabric_pd_active_i9                                      => fabric_pd_active_i(8)
       , fabric_pd_active_i10                                     => fabric_pd_active_i(9)
       , fabric_pd_active_i11                                     => fabric_pd_active_i(10)
       , fabric_pd_active_i12                                     => fabric_pd_active_i(11)
       , fabric_pd_active_i13                                     => fabric_pd_active_i(12)
       , fabric_pd_active_i14                                     => fabric_pd_active_i(13)
       , fabric_pd_active_i15                                     => fabric_pd_active_i(14)
       , fabric_pd_active_i16                                     => fabric_pd_active_i(15)
       , fabric_pd_active_i17                                     => fabric_pd_active_i(16)
       , fabric_pd_active_i18                                     => fabric_pd_active_i(17)
       , fabric_pd_active_i19                                     => fabric_pd_active_i(18)
       , fabric_pd_active_i20                                     => fabric_pd_active_i(19)
       , fabric_pd_active_i21                                     => fabric_pd_active_i(20)
       , fabric_pd_active_i22                                     => fabric_pd_active_i(21)
       , fabric_pd_active_i23                                     => fabric_pd_active_i(22)
       , fabric_pd_active_i24                                     => fabric_pd_active_i(23)
       , fabric_otp_user_suppadd_i                                => fabric_otp_user_suppadd_i
       , fabric_mrepair_fuse_pdn_i                                => fabric_mrepair_fuse_pdn_i
       , fabric_otp_security_scanin_i1                            => fabric_otp_security_scanin_i(0)
       , fabric_otp_security_scanin_i2                            => fabric_otp_security_scanin_i(1)
       , fabric_otp_security_scanin_i3                            => fabric_otp_security_scanin_i(2)
       , fabric_otp_security_scanin_i4                            => fabric_otp_security_scanin_i(3)
       , fabric_otp_security_scanin_i5                            => fabric_otp_security_scanin_i(4)
       , fabric_end_encoding_i                                    => fabric_end_encoding_i
       , fabric_jtag_tdo_usr2_i                                   => fabric_jtag_tdo_usr2_i
       , fabric_mrepair_fuse_wordlock_i                           => fabric_mrepair_fuse_wordlock_i
       , fabric_otp_user_prgwidth_i1                              => fabric_otp_user_prgwidth_i(0)
       , fabric_otp_user_prgwidth_i2                              => fabric_otp_user_prgwidth_i(1)
       , fabric_otp_user_prgwidth_i3                              => fabric_otp_user_prgwidth_i(2)
       , fabric_otp_user_read_i                                   => fabric_otp_user_read_i
       , fabric_mrepair_fuse_add_i1                               => fabric_mrepair_fuse_add_i(0)
       , fabric_mrepair_fuse_add_i2                               => fabric_mrepair_fuse_add_i(1)
       , fabric_mrepair_fuse_add_i3                               => fabric_mrepair_fuse_add_i(2)
       , fabric_mrepair_fuse_add_i4                               => fabric_mrepair_fuse_add_i(3)
       , fabric_mrepair_fuse_add_i5                               => fabric_mrepair_fuse_add_i(4)
       , fabric_mrepair_fuse_add_i6                               => fabric_mrepair_fuse_add_i(5)
       , fabric_mrepair_fuse_add_i7                               => fabric_mrepair_fuse_add_i(6)
       , fabric_mrepair_fuse_bistmode_i                           => fabric_mrepair_fuse_bistmode_i
       , fabric_jtag_tdo_usr1_i                                   => fabric_jtag_tdo_usr1_i
       , fabric_otp_cfg_clk_fab_en_i                              => fabric_otp_cfg_clk_fab_en_i
       , fabric_io_in_i1                                          => fabric_io_in_i(0)
       , fabric_io_in_i2                                          => fabric_io_in_i(1)
       , fabric_io_in_i3                                          => fabric_io_in_i(2)
       , fabric_io_in_i4                                          => fabric_io_in_i(3)
       , fabric_io_in_i5                                          => fabric_io_in_i(4)
       , fabric_io_in_i6                                          => fabric_io_in_i(5)
       , fabric_io_in_i7                                          => fabric_io_in_i(6)
       , fabric_io_in_i8                                          => fabric_io_in_i(7)
       , fabric_io_in_i9                                          => fabric_io_in_i(8)
       , fabric_io_in_i10                                         => fabric_io_in_i(9)
       , fabric_io_in_i11                                         => fabric_io_in_i(10)
       , fabric_io_in_i12                                         => fabric_io_in_i(11)
       , fabric_io_in_i13                                         => fabric_io_in_i(12)
       , fabric_io_in_i14                                         => fabric_io_in_i(13)
       , fabric_io_in_i15                                         => fabric_io_in_i(14)
       , fabric_io_in_i16                                         => fabric_io_in_i(15)
       , fabric_io_in_i17                                         => fabric_io_in_i(16)
       , fabric_io_in_i18                                         => fabric_io_in_i(17)
       , fabric_io_in_i19                                         => fabric_io_in_i(18)
       , fabric_io_in_i20                                         => fabric_io_in_i(19)
       , fabric_io_in_i21                                         => fabric_io_in_i(20)
       , fabric_io_in_i22                                         => fabric_io_in_i(21)
       , fabric_io_in_i23                                         => fabric_io_in_i(22)
       , fabric_io_in_i24                                         => fabric_io_in_i(23)
       , fabric_io_in_i25                                         => fabric_io_in_i(24)
       , fabric_sif_load_en_i1                                    => fabric_sif_load_en_i(0)
       , fabric_sif_load_en_i2                                    => fabric_sif_load_en_i(1)
       , fabric_sif_load_en_i3                                    => fabric_sif_load_en_i(2)
       , fabric_sif_load_en_i4                                    => fabric_sif_load_en_i(3)
       , fabric_sif_load_en_i5                                    => fabric_sif_load_en_i(4)
       , fabric_sif_load_en_i6                                    => fabric_sif_load_en_i(5)
       , fabric_sif_load_en_i7                                    => fabric_sif_load_en_i(6)
       , fabric_sif_load_en_i8                                    => fabric_sif_load_en_i(7)
       , fabric_sif_load_en_i9                                    => fabric_sif_load_en_i(8)
       , fabric_sif_load_en_i10                                   => fabric_sif_load_en_i(9)
       , fabric_sif_load_en_i11                                   => fabric_sif_load_en_i(10)
       , fabric_sif_load_en_i12                                   => fabric_sif_load_en_i(11)
       , fabric_sif_load_en_i13                                   => fabric_sif_load_en_i(12)
       , fabric_sif_load_en_i14                                   => fabric_sif_load_en_i(13)
       , fabric_sif_load_en_i15                                   => fabric_sif_load_en_i(14)
       , fabric_sif_load_en_i16                                   => fabric_sif_load_en_i(15)
       , fabric_sif_load_en_i17                                   => fabric_sif_load_en_i(16)
       , fabric_sif_load_en_i18                                   => fabric_sif_load_en_i(17)
       , fabric_sif_load_en_i19                                   => fabric_sif_load_en_i(18)
       , fabric_sif_load_en_i20                                   => fabric_sif_load_en_i(19)
       , fabric_sif_load_en_i21                                   => fabric_sif_load_en_i(20)
       , fabric_sif_load_en_i22                                   => fabric_sif_load_en_i(21)
       , fabric_sif_load_en_i23                                   => fabric_sif_load_en_i(22)
       , fabric_sif_load_en_i24                                   => fabric_sif_load_en_i(23)
       , fabric_mrepair_fuse_din_i1                               => fabric_mrepair_fuse_din_i(0)
       , fabric_mrepair_fuse_din_i2                               => fabric_mrepair_fuse_din_i(1)
       , fabric_mrepair_fuse_din_i3                               => fabric_mrepair_fuse_din_i(2)
       , fabric_mrepair_fuse_din_i4                               => fabric_mrepair_fuse_din_i(3)
       , fabric_mrepair_fuse_din_i5                               => fabric_mrepair_fuse_din_i(4)
       , fabric_mrepair_fuse_din_i6                               => fabric_mrepair_fuse_din_i(5)
       , fabric_mrepair_fuse_din_i7                               => fabric_mrepair_fuse_din_i(6)
       , fabric_mrepair_fuse_din_i8                               => fabric_mrepair_fuse_din_i(7)
       , fabric_mrepair_fuse_din_i9                               => fabric_mrepair_fuse_din_i(8)
       , fabric_mrepair_fuse_din_i10                              => fabric_mrepair_fuse_din_i(9)
       , fabric_mrepair_fuse_din_i11                              => fabric_mrepair_fuse_din_i(10)
       , fabric_mrepair_fuse_din_i12                              => fabric_mrepair_fuse_din_i(11)
       , fabric_mrepair_fuse_din_i13                              => fabric_mrepair_fuse_din_i(12)
       , fabric_mrepair_fuse_din_i14                              => fabric_mrepair_fuse_din_i(13)
       , fabric_mrepair_fuse_din_i15                              => fabric_mrepair_fuse_din_i(14)
       , fabric_mrepair_fuse_din_i16                              => fabric_mrepair_fuse_din_i(15)
       , fabric_mrepair_fuse_din_i17                              => fabric_mrepair_fuse_din_i(16)
       , fabric_mrepair_fuse_din_i18                              => fabric_mrepair_fuse_din_i(17)
       , fabric_mrepair_fuse_din_i19                              => fabric_mrepair_fuse_din_i(18)
       , fabric_mrepair_fuse_din_i20                              => fabric_mrepair_fuse_din_i(19)
       , fabric_mrepair_fuse_din_i21                              => fabric_mrepair_fuse_din_i(20)
       , fabric_mrepair_fuse_din_i22                              => fabric_mrepair_fuse_din_i(21)
       , fabric_mrepair_fuse_din_i23                              => fabric_mrepair_fuse_din_i(22)
       , fabric_mrepair_fuse_din_i24                              => fabric_mrepair_fuse_din_i(23)
       , fabric_mrepair_fuse_din_i25                              => fabric_mrepair_fuse_din_i(24)
       , fabric_mrepair_fuse_din_i26                              => fabric_mrepair_fuse_din_i(25)
       , fabric_mrepair_fuse_din_i27                              => fabric_mrepair_fuse_din_i(26)
       , fabric_mrepair_fuse_din_i28                              => fabric_mrepair_fuse_din_i(27)
       , fabric_mrepair_fuse_din_i29                              => fabric_mrepair_fuse_din_i(28)
       , fabric_mrepair_fuse_din_i30                              => fabric_mrepair_fuse_din_i(29)
       , fabric_mrepair_fuse_din_i31                              => fabric_mrepair_fuse_din_i(30)
       , fabric_mrepair_fuse_din_i32                              => fabric_mrepair_fuse_din_i(31)
       , fabric_mrepair_fuse_din_i33                              => fabric_mrepair_fuse_din_i(32)
       , fabric_mrepair_fuse_din_i34                              => fabric_mrepair_fuse_din_i(33)
       , fabric_mrepair_fuse_din_i35                              => fabric_mrepair_fuse_din_i(34)
       , fabric_mrepair_fuse_din_i36                              => fabric_mrepair_fuse_din_i(35)
       , fabric_mrepair_fuse_din_i37                              => fabric_mrepair_fuse_din_i(36)
       , fabric_mrepair_fuse_din_i38                              => fabric_mrepair_fuse_din_i(37)
       , fabric_mrepair_fuse_din_i39                              => fabric_mrepair_fuse_din_i(38)
       , fabric_otp_apb_addr_i1                                   => fabric_otp_apb_addr_i(0)
       , fabric_otp_apb_addr_i2                                   => fabric_otp_apb_addr_i(1)
       , fabric_otp_apb_addr_i3                                   => fabric_otp_apb_addr_i(2)
       , fabric_otp_apb_addr_i4                                   => fabric_otp_apb_addr_i(3)
       , fabric_otp_apb_addr_i5                                   => fabric_otp_apb_addr_i(4)
       , fabric_otp_apb_addr_i6                                   => fabric_otp_apb_addr_i(5)
       , fabric_otp_apb_addr_i7                                   => fabric_otp_apb_addr_i(6)
       , fabric_otp_apb_addr_i8                                   => fabric_otp_apb_addr_i(7)
       , fabric_otp_apb_addr_i9                                   => fabric_otp_apb_addr_i(8)
       , fabric_otp_apb_addr_i10                                  => fabric_otp_apb_addr_i(9)
       , fabric_otp_apb_addr_i11                                  => fabric_otp_apb_addr_i(10)
       , fabric_otp_apb_addr_i12                                  => fabric_otp_apb_addr_i(11)
       , fabric_otp_apb_addr_i13                                  => fabric_otp_apb_addr_i(12)
       , fabric_otp_apb_addr_i14                                  => fabric_otp_apb_addr_i(13)
       , fabric_otp_apb_addr_i15                                  => fabric_otp_apb_addr_i(14)
       , fabric_otp_apb_addr_i16                                  => fabric_otp_apb_addr_i(15)
       , fabric_otp_apb_addr_i17                                  => fabric_otp_apb_addr_i(16)
       , fabric_otp_apb_addr_i18                                  => fabric_otp_apb_addr_i(17)
       , fabric_otp_apb_addr_i19                                  => fabric_otp_apb_addr_i(18)
       , fabric_otp_apb_addr_i20                                  => fabric_otp_apb_addr_i(19)
       , fabric_otp_apb_addr_i21                                  => fabric_otp_apb_addr_i(20)
       , fabric_otp_apb_addr_i22                                  => fabric_otp_apb_addr_i(21)
       , fabric_otp_apb_addr_i23                                  => fabric_otp_apb_addr_i(22)
       , fabric_otp_apb_addr_i24                                  => fabric_otp_apb_addr_i(23)
       , fabric_otp_apb_addr_i25                                  => fabric_otp_apb_addr_i(24)
       , fabric_otp_apb_addr_i26                                  => fabric_otp_apb_addr_i(25)
       , fabric_otp_apb_addr_i27                                  => fabric_otp_apb_addr_i(26)
       , fabric_otp_apb_addr_i28                                  => fabric_otp_apb_addr_i(27)
       , fabric_otp_apb_addr_i29                                  => fabric_otp_apb_addr_i(28)
       , fabric_otp_apb_addr_i30                                  => fabric_otp_apb_addr_i(29)
       , fabric_otp_apb_addr_i31                                  => fabric_otp_apb_addr_i(30)
       , fabric_otp_apb_addr_i32                                  => fabric_otp_apb_addr_i(31)
       , fabric_otp_apb_sel_i                                     => fabric_otp_apb_sel_i
       , fabric_mrepair_fuse_rbact1_i                             => fabric_mrepair_fuse_rbact1_i
       , fabric_mrepair_fuse_configreg_i1                         => fabric_mrepair_fuse_configreg_i(0)
       , fabric_mrepair_fuse_configreg_i2                         => fabric_mrepair_fuse_configreg_i(1)
       , fabric_mrepair_fuse_configreg_i3                         => fabric_mrepair_fuse_configreg_i(2)
       , fabric_mrepair_fuse_configreg_i4                         => fabric_mrepair_fuse_configreg_i(3)
       , fabric_mrepair_fuse_configreg_i5                         => fabric_mrepair_fuse_configreg_i(4)
       , fabric_mrepair_fuse_configreg_i6                         => fabric_mrepair_fuse_configreg_i(5)
       , fabric_mrepair_fuse_configreg_i7                         => fabric_mrepair_fuse_configreg_i(6)
       , fabric_mrepair_fuse_configreg_i8                         => fabric_mrepair_fuse_configreg_i(7)
       , fabric_mrepair_fuse_configreg_i9                         => fabric_mrepair_fuse_configreg_i(8)
       , fabric_mrepair_fuse_configreg_i10                        => fabric_mrepair_fuse_configreg_i(9)
       , fabric_mrepair_fuse_configreg_i11                        => fabric_mrepair_fuse_configreg_i(10)
       , fabric_mrepair_fuse_configreg_i12                        => fabric_mrepair_fuse_configreg_i(11)
       , fabric_mrepair_fuse_configreg_i13                        => fabric_mrepair_fuse_configreg_i(12)
       , fabric_mrepair_fuse_configreg_i14                        => fabric_mrepair_fuse_configreg_i(13)
       , fabric_mrepair_fuse_configreg_i15                        => fabric_mrepair_fuse_configreg_i(14)
       , fabric_mrepair_fuse_configreg_i16                        => fabric_mrepair_fuse_configreg_i(15)
       , fabric_mrepair_fuse_configreg_i17                        => fabric_mrepair_fuse_configreg_i(16)
       , fabric_mrepair_fuse_configreg_i18                        => fabric_mrepair_fuse_configreg_i(17)
       , fabric_mrepair_fuse_configreg_i19                        => fabric_mrepair_fuse_configreg_i(18)
       , fabric_mrepair_fuse_configreg_i20                        => fabric_mrepair_fuse_configreg_i(19)
       , fabric_mrepair_fuse_configreg_i21                        => fabric_mrepair_fuse_configreg_i(20)
       , fabric_mrepair_fuse_configreg_i22                        => fabric_mrepair_fuse_configreg_i(21)
       , fabric_mrepair_fuse_configreg_i23                        => fabric_mrepair_fuse_configreg_i(22)
       , fabric_mrepair_fuse_configreg_i24                        => fabric_mrepair_fuse_configreg_i(23)
       , fabric_mrepair_fuse_configreg_i25                        => fabric_mrepair_fuse_configreg_i(24)
       , fabric_mrepair_fuse_configreg_i26                        => fabric_mrepair_fuse_configreg_i(25)
       , fabric_mrepair_fuse_configreg_i27                        => fabric_mrepair_fuse_configreg_i(26)
       , fabric_mrepair_fuse_configreg_i28                        => fabric_mrepair_fuse_configreg_i(27)
       , fabric_mrepair_fuse_configreg_i29                        => fabric_mrepair_fuse_configreg_i(28)
       , fabric_mrepair_fuse_configreg_i30                        => fabric_mrepair_fuse_configreg_i(29)
       , fabric_mrepair_fuse_configreg_i31                        => fabric_mrepair_fuse_configreg_i(30)
       , fabric_mrepair_fuse_configreg_i32                        => fabric_mrepair_fuse_configreg_i(31)
       , fabric_otp_cfg_fabric_apb_en_i                           => fabric_otp_cfg_fabric_apb_en_i
       , fabric_data_shift_en_i                                   => fabric_data_shift_en_i
       , fabric_lowskew_i21                                       => fabric_lowskew_i21
       , fabric_direct_data_i1                                    => fabric_direct_data_i(0)
       , fabric_direct_data_i2                                    => fabric_direct_data_i(1)
       , fabric_direct_data_i3                                    => fabric_direct_data_i(2)
       , fabric_direct_data_i4                                    => fabric_direct_data_i(3)
       , fabric_direct_data_i5                                    => fabric_direct_data_i(4)
       , fabric_direct_data_i6                                    => fabric_direct_data_i(5)
       , fabric_direct_data_i7                                    => fabric_direct_data_i(6)
       , fabric_direct_data_i8                                    => fabric_direct_data_i(7)
       , fabric_direct_data_i9                                    => fabric_direct_data_i(8)
       , fabric_direct_data_i10                                   => fabric_direct_data_i(9)
       , fabric_direct_data_i11                                   => fabric_direct_data_i(10)
       , fabric_direct_data_i12                                   => fabric_direct_data_i(11)
       , fabric_direct_data_i13                                   => fabric_direct_data_i(12)
       , fabric_direct_data_i14                                   => fabric_direct_data_i(13)
       , fabric_direct_data_i15                                   => fabric_direct_data_i(14)
       , fabric_direct_data_i16                                   => fabric_direct_data_i(15)
       , fabric_direct_data_i17                                   => fabric_direct_data_i(16)
       , fabric_direct_data_i18                                   => fabric_direct_data_i(17)
       , fabric_direct_data_i19                                   => fabric_direct_data_i(18)
       , fabric_direct_data_i20                                   => fabric_direct_data_i(19)
       , fabric_direct_data_i21                                   => fabric_direct_data_i(20)
       , fabric_direct_data_i22                                   => fabric_direct_data_i(21)
       , fabric_direct_data_i23                                   => fabric_direct_data_i(22)
       , fabric_direct_data_i24                                   => fabric_direct_data_i(23)
       , fabric_direct_data_i25                                   => fabric_direct_data_i(24)
       , fabric_direct_data_i26                                   => fabric_direct_data_i(25)
       , fabric_direct_data_i27                                   => fabric_direct_data_i(26)
       , fabric_direct_data_i28                                   => fabric_direct_data_i(27)
       , fabric_direct_data_i29                                   => fabric_direct_data_i(28)
       , fabric_direct_data_i30                                   => fabric_direct_data_i(29)
       , fabric_direct_data_i31                                   => fabric_direct_data_i(30)
       , fabric_direct_data_i32                                   => fabric_direct_data_i(31)
       , fabric_otp_user_pdn_i                                    => fabric_otp_user_pdn_i
       , fabric_io_oe_i1                                          => fabric_io_oe_i(0)
       , fabric_io_oe_i2                                          => fabric_io_oe_i(1)
       , fabric_io_oe_i3                                          => fabric_io_oe_i(2)
       , fabric_io_oe_i4                                          => fabric_io_oe_i(3)
       , fabric_io_oe_i5                                          => fabric_io_oe_i(4)
       , fabric_io_oe_i6                                          => fabric_io_oe_i(5)
       , fabric_io_oe_i7                                          => fabric_io_oe_i(6)
       , fabric_io_oe_i8                                          => fabric_io_oe_i(7)
       , fabric_io_oe_i9                                          => fabric_io_oe_i(8)
       , fabric_io_oe_i10                                         => fabric_io_oe_i(9)
       , fabric_io_oe_i11                                         => fabric_io_oe_i(10)
       , fabric_io_oe_i12                                         => fabric_io_oe_i(11)
       , fabric_io_oe_i13                                         => fabric_io_oe_i(12)
       , fabric_io_oe_i14                                         => fabric_io_oe_i(13)
       , fabric_io_oe_i15                                         => fabric_io_oe_i(14)
       , fabric_io_oe_i16                                         => fabric_io_oe_i(15)
       , fabric_io_oe_i17                                         => fabric_io_oe_i(16)
       , fabric_io_oe_i18                                         => fabric_io_oe_i(17)
       , fabric_io_oe_i19                                         => fabric_io_oe_i(18)
       , fabric_io_oe_i20                                         => fabric_io_oe_i(19)
       , fabric_io_oe_i21                                         => fabric_io_oe_i(20)
       , fabric_io_oe_i22                                         => fabric_io_oe_i(21)
       , fabric_io_oe_i23                                         => fabric_io_oe_i(22)
       , fabric_io_oe_i24                                         => fabric_io_oe_i(23)
       , fabric_io_oe_i25                                         => fabric_io_oe_i(24)
       , fabric_parusr_data_i1                                    => fabric_parusr_data_i(0)
       , fabric_parusr_data_i2                                    => fabric_parusr_data_i(1)
       , fabric_parusr_data_i3                                    => fabric_parusr_data_i(2)
       , fabric_parusr_data_i4                                    => fabric_parusr_data_i(3)
       , fabric_parusr_data_i5                                    => fabric_parusr_data_i(4)
       , fabric_parusr_data_i6                                    => fabric_parusr_data_i(5)
       , fabric_parusr_data_i7                                    => fabric_parusr_data_i(6)
       , fabric_parusr_data_i8                                    => fabric_parusr_data_i(7)
       , fabric_parusr_data_i9                                    => fabric_parusr_data_i(8)
       , fabric_parusr_data_i10                                   => fabric_parusr_data_i(9)
       , fabric_parusr_data_i11                                   => fabric_parusr_data_i(10)
       , fabric_parusr_data_i12                                   => fabric_parusr_data_i(11)
       , fabric_parusr_data_i13                                   => fabric_parusr_data_i(12)
       , fabric_parusr_data_i14                                   => fabric_parusr_data_i(13)
       , fabric_parusr_data_i15                                   => fabric_parusr_data_i(14)
       , fabric_parusr_data_i16                                   => fabric_parusr_data_i(15)
       , fabric_otp_apb_write_i                                   => fabric_otp_apb_write_i
       , fabric_otp_security_testmode_i                           => fabric_otp_security_testmode_i
       , fabric_system_data_to_mem_bist_i1                        => fabric_system_data_to_mem_bist_i(0)
       , fabric_system_data_to_mem_bist_i2                        => fabric_system_data_to_mem_bist_i(1)
       , fabric_system_data_to_mem_bist_i3                        => fabric_system_data_to_mem_bist_i(2)
       , fabric_system_data_to_mem_bist_i4                        => fabric_system_data_to_mem_bist_i(3)
       , fabric_system_data_to_mem_bist_i5                        => fabric_system_data_to_mem_bist_i(4)
       , fabric_system_data_to_mem_bist_i6                        => fabric_system_data_to_mem_bist_i(5)
       , fabric_system_data_to_mem_bist_i7                        => fabric_system_data_to_mem_bist_i(6)
       , fabric_system_data_to_mem_bist_i8                        => fabric_system_data_to_mem_bist_i(7)
       , fabric_system_data_to_mem_bist_i9                        => fabric_system_data_to_mem_bist_i(8)
       , fabric_system_data_to_mem_bist_i10                       => fabric_system_data_to_mem_bist_i(9)
       , fabric_system_data_to_mem_bist_i11                       => fabric_system_data_to_mem_bist_i(10)
       , fabric_system_data_to_mem_bist_i12                       => fabric_system_data_to_mem_bist_i(11)
       , fabric_system_data_to_mem_bist_i13                       => fabric_system_data_to_mem_bist_i(12)
       , fabric_system_data_to_mem_bist_i14                       => fabric_system_data_to_mem_bist_i(13)
       , fabric_system_data_to_mem_bist_i15                       => fabric_system_data_to_mem_bist_i(14)
       , fabric_system_data_to_mem_bist_i16                       => fabric_system_data_to_mem_bist_i(15)
       , fabric_system_data_to_mem_bist_i17                       => fabric_system_data_to_mem_bist_i(16)
       , fabric_system_data_to_mem_bist_i18                       => fabric_system_data_to_mem_bist_i(17)
       , fabric_system_data_to_mem_bist_i19                       => fabric_system_data_to_mem_bist_i(18)
       , fabric_system_data_to_mem_bist_i20                       => fabric_system_data_to_mem_bist_i(19)
       , fabric_system_data_to_mem_bist_i21                       => fabric_system_data_to_mem_bist_i(20)
       , fabric_system_data_to_mem_bist_i22                       => fabric_system_data_to_mem_bist_i(21)
       , fabric_system_data_to_mem_bist_i23                       => fabric_system_data_to_mem_bist_i(22)
       , fabric_system_data_to_mem_bist_i24                       => fabric_system_data_to_mem_bist_i(23)
       , fabric_tst_atpg_mrepair_i                                => fabric_tst_atpg_mrepair_i
       , fabric_mrepair_fuse_tstscanenable_i                      => fabric_mrepair_fuse_tstscanenable_i
       , fabric_otp_security_bistmode_i                           => fabric_otp_security_bistmode_i
       , fabric_lowskew_i22                                       => fabric_lowskew_i22
       , fabric_lowskew_i23                                       => fabric_lowskew_i23
       , fabric_lowskew_i20                                       => fabric_lowskew_i20
       , fabric_otp_user_configreg_i1                             => fabric_otp_user_configreg_i(0)
       , fabric_otp_user_configreg_i2                             => fabric_otp_user_configreg_i(1)
       , fabric_otp_user_configreg_i3                             => fabric_otp_user_configreg_i(2)
       , fabric_otp_user_configreg_i4                             => fabric_otp_user_configreg_i(3)
       , fabric_otp_user_configreg_i5                             => fabric_otp_user_configreg_i(4)
       , fabric_otp_user_configreg_i6                             => fabric_otp_user_configreg_i(5)
       , fabric_otp_user_configreg_i7                             => fabric_otp_user_configreg_i(6)
       , fabric_otp_user_configreg_i8                             => fabric_otp_user_configreg_i(7)
       , fabric_otp_user_configreg_i9                             => fabric_otp_user_configreg_i(8)
       , fabric_otp_user_configreg_i10                            => fabric_otp_user_configreg_i(9)
       , fabric_otp_user_configreg_i11                            => fabric_otp_user_configreg_i(10)
       , fabric_otp_user_configreg_i12                            => fabric_otp_user_configreg_i(11)
       , fabric_otp_user_configreg_i13                            => fabric_otp_user_configreg_i(12)
       , fabric_otp_user_configreg_i14                            => fabric_otp_user_configreg_i(13)
       , fabric_otp_user_configreg_i15                            => fabric_otp_user_configreg_i(14)
       , fabric_otp_user_configreg_i16                            => fabric_otp_user_configreg_i(15)
       , fabric_otp_user_configreg_i17                            => fabric_otp_user_configreg_i(16)
       , fabric_otp_user_configreg_i18                            => fabric_otp_user_configreg_i(17)
       , fabric_otp_user_configreg_i19                            => fabric_otp_user_configreg_i(18)
       , fabric_otp_user_configreg_i20                            => fabric_otp_user_configreg_i(19)
       , fabric_otp_user_configreg_i21                            => fabric_otp_user_configreg_i(20)
       , fabric_otp_user_configreg_i22                            => fabric_otp_user_configreg_i(21)
       , fabric_otp_user_configreg_i23                            => fabric_otp_user_configreg_i(22)
       , fabric_otp_user_configreg_i24                            => fabric_otp_user_configreg_i(23)
       , fabric_otp_user_configreg_i25                            => fabric_otp_user_configreg_i(24)
       , fabric_otp_user_configreg_i26                            => fabric_otp_user_configreg_i(25)
       , fabric_otp_user_configreg_i27                            => fabric_otp_user_configreg_i(26)
       , fabric_otp_user_configreg_i28                            => fabric_otp_user_configreg_i(27)
       , fabric_otp_user_configreg_i29                            => fabric_otp_user_configreg_i(28)
       , fabric_otp_user_configreg_i30                            => fabric_otp_user_configreg_i(29)
       , fabric_otp_user_configreg_i31                            => fabric_otp_user_configreg_i(30)
       , fabric_otp_user_configreg_i32                            => fabric_otp_user_configreg_i(31)
       , fabric_otp_user_tst_scanin_i1                            => fabric_otp_user_tst_scanin_i(0)
       , fabric_otp_user_tst_scanin_i2                            => fabric_otp_user_tst_scanin_i(1)
       , fabric_otp_user_tst_scanin_i3                            => fabric_otp_user_tst_scanin_i(2)
       , fabric_otp_user_tst_scanin_i4                            => fabric_otp_user_tst_scanin_i(3)
       , fabric_otp_user_tst_scanin_i5                            => fabric_otp_user_tst_scanin_i(4)
       , fabric_sif_update_en_i1                                  => fabric_sif_update_en_i(0)
       , fabric_sif_update_en_i2                                  => fabric_sif_update_en_i(1)
       , fabric_sif_update_en_i3                                  => fabric_sif_update_en_i(2)
       , fabric_sif_update_en_i4                                  => fabric_sif_update_en_i(3)
       , fabric_sif_update_en_i5                                  => fabric_sif_update_en_i(4)
       , fabric_sif_update_en_i6                                  => fabric_sif_update_en_i(5)
       , fabric_sif_update_en_i7                                  => fabric_sif_update_en_i(6)
       , fabric_sif_update_en_i8                                  => fabric_sif_update_en_i(7)
       , fabric_sif_update_en_i9                                  => fabric_sif_update_en_i(8)
       , fabric_sif_update_en_i10                                 => fabric_sif_update_en_i(9)
       , fabric_sif_update_en_i11                                 => fabric_sif_update_en_i(10)
       , fabric_sif_update_en_i12                                 => fabric_sif_update_en_i(11)
       , fabric_sif_update_en_i13                                 => fabric_sif_update_en_i(12)
       , fabric_sif_update_en_i14                                 => fabric_sif_update_en_i(13)
       , fabric_sif_update_en_i15                                 => fabric_sif_update_en_i(14)
       , fabric_sif_update_en_i16                                 => fabric_sif_update_en_i(15)
       , fabric_sif_update_en_i17                                 => fabric_sif_update_en_i(16)
       , fabric_sif_update_en_i18                                 => fabric_sif_update_en_i(17)
       , fabric_sif_update_en_i19                                 => fabric_sif_update_en_i(18)
       , fabric_sif_update_en_i20                                 => fabric_sif_update_en_i(19)
       , fabric_sif_update_en_i21                                 => fabric_sif_update_en_i(20)
       , fabric_sif_update_en_i22                                 => fabric_sif_update_en_i(21)
       , fabric_sif_update_en_i23                                 => fabric_sif_update_en_i(22)
       , fabric_sif_update_en_i24                                 => fabric_sif_update_en_i(23)
       , fabric_mrepair_por_i                                     => fabric_mrepair_por_i
       , fabric_mrepair_rst_n_i                                   => fabric_mrepair_rst_n_i
       , fabric_mrepair_initn_i                                   => fabric_mrepair_initn_i
       , fabric_spare_i1                                          => fabric_spare_i(0)
       , fabric_spare_i2                                          => fabric_spare_i(1)
       , fabric_spare_i3                                          => fabric_spare_i(2)
       , fabric_mrepair_fuse_bbad_o                               => fabric_mrepair_fuse_bbad_o
       , fabric_jtag_trst_n_o                                     => fabric_jtag_trst_n_o
       , fabric_debug_direct_permission_write_o1                  => fabric_debug_direct_permission_write_o(0)
       , fabric_debug_direct_permission_write_o2                  => fabric_debug_direct_permission_write_o(1)
       , fabric_debug_direct_permission_write_o3                  => fabric_debug_direct_permission_write_o(2)
       , fabric_debug_direct_permission_write_o4                  => fabric_debug_direct_permission_write_o(3)
       , fabric_otp_security_bist_end1_o                          => fabric_otp_security_bist_end1_o
       , fabric_parusr_data_val_o                                 => fabric_parusr_data_val_o
       , fabric_debug_lock_reg_o                                  => fabric_debug_lock_reg_o
       , fabric_debug_security_error_read_o                       => fabric_debug_security_error_read_o
       , fabric_mrepair_fuse_tstscanout_o1                        => fabric_mrepair_fuse_tstscanout_o(0)
       , fabric_mrepair_fuse_tstscanout_o2                        => fabric_mrepair_fuse_tstscanout_o(1)
       , fabric_mrepair_fuse_tstscanout_o3                        => fabric_mrepair_fuse_tstscanout_o(2)
       , fabric_mrepair_fuse_tstscanout_o4                        => fabric_mrepair_fuse_tstscanout_o(3)
       , fabric_mrepair_fuse_tstscanout_o5                        => fabric_mrepair_fuse_tstscanout_o(4)
       , fabric_otp_user_tst_scanout_o1                           => fabric_otp_user_tst_scanout_o(0)
       , fabric_otp_user_tst_scanout_o2                           => fabric_otp_user_tst_scanout_o(1)
       , fabric_otp_user_tst_scanout_o3                           => fabric_otp_user_tst_scanout_o(2)
       , fabric_otp_user_tst_scanout_o4                           => fabric_otp_user_tst_scanout_o(3)
       , fabric_otp_user_tst_scanout_o5                           => fabric_otp_user_tst_scanout_o(4)
       , fabric_sif_update_en_to_bist_o1                          => fabric_sif_update_en_to_bist_o(0)
       , fabric_sif_update_en_to_bist_o2                          => fabric_sif_update_en_to_bist_o(1)
       , fabric_sif_update_en_to_bist_o3                          => fabric_sif_update_en_to_bist_o(2)
       , fabric_sif_update_en_to_bist_o4                          => fabric_sif_update_en_to_bist_o(3)
       , fabric_sif_update_en_to_bist_o5                          => fabric_sif_update_en_to_bist_o(4)
       , fabric_sif_update_en_to_bist_o6                          => fabric_sif_update_en_to_bist_o(5)
       , fabric_sif_update_en_to_bist_o7                          => fabric_sif_update_en_to_bist_o(6)
       , fabric_sif_update_en_to_bist_o8                          => fabric_sif_update_en_to_bist_o(7)
       , fabric_sif_update_en_to_bist_o9                          => fabric_sif_update_en_to_bist_o(8)
       , fabric_sif_update_en_to_bist_o10                         => fabric_sif_update_en_to_bist_o(9)
       , fabric_sif_update_en_to_bist_o11                         => fabric_sif_update_en_to_bist_o(10)
       , fabric_sif_update_en_to_bist_o12                         => fabric_sif_update_en_to_bist_o(11)
       , fabric_sif_update_en_to_bist_o13                         => fabric_sif_update_en_to_bist_o(12)
       , fabric_sif_update_en_to_bist_o14                         => fabric_sif_update_en_to_bist_o(13)
       , fabric_sif_update_en_to_bist_o15                         => fabric_sif_update_en_to_bist_o(14)
       , fabric_sif_update_en_to_bist_o16                         => fabric_sif_update_en_to_bist_o(15)
       , fabric_sif_update_en_to_bist_o17                         => fabric_sif_update_en_to_bist_o(16)
       , fabric_sif_update_en_to_bist_o18                         => fabric_sif_update_en_to_bist_o(17)
       , fabric_sif_update_en_to_bist_o19                         => fabric_sif_update_en_to_bist_o(18)
       , fabric_sif_update_en_to_bist_o20                         => fabric_sif_update_en_to_bist_o(19)
       , fabric_sif_update_en_to_bist_o21                         => fabric_sif_update_en_to_bist_o(20)
       , fabric_sif_update_en_to_bist_o22                         => fabric_sif_update_en_to_bist_o(21)
       , fabric_sif_update_en_to_bist_o23                         => fabric_sif_update_en_to_bist_o(22)
       , fabric_sif_update_en_to_bist_o24                         => fabric_sif_update_en_to_bist_o(23)
       , fabric_otp_user_locked_o                                 => fabric_otp_user_locked_o
       , fabric_otp_security_bist_bad_o                           => fabric_otp_security_bist_bad_o
       , fabric_debug_frame_permission_frame_o1                   => fabric_debug_frame_permission_frame_o(0)
       , fabric_debug_frame_permission_frame_o2                   => fabric_debug_frame_permission_frame_o(1)
       , fabric_debug_frame_permission_frame_o3                   => fabric_debug_frame_permission_frame_o(2)
       , fabric_debug_frame_permission_frame_o4                   => fabric_debug_frame_permission_frame_o(3)
       , fabric_otp_user_pwok_o                                   => fabric_otp_user_pwok_o
       , fabric_otp_user_bend2_o                                  => fabric_otp_user_bend2_o
       , fabric_mrepair_fuse_ded_o                                => fabric_mrepair_fuse_ded_o
       , fabric_debug_access_reg_data_ready_o                     => fabric_debug_access_reg_data_ready_o
       , fabric_data_to_bist_o1                                   => fabric_data_to_bist_o(0)
       , fabric_data_to_bist_o2                                   => fabric_data_to_bist_o(1)
       , fabric_data_to_bist_o3                                   => fabric_data_to_bist_o(2)
       , fabric_data_to_bist_o4                                   => fabric_data_to_bist_o(3)
       , fabric_data_to_bist_o5                                   => fabric_data_to_bist_o(4)
       , fabric_data_to_bist_o6                                   => fabric_data_to_bist_o(5)
       , fabric_data_to_bist_o7                                   => fabric_data_to_bist_o(6)
       , fabric_data_to_bist_o8                                   => fabric_data_to_bist_o(7)
       , fabric_data_to_bist_o9                                   => fabric_data_to_bist_o(8)
       , fabric_data_to_bist_o10                                  => fabric_data_to_bist_o(9)
       , fabric_data_to_bist_o11                                  => fabric_data_to_bist_o(10)
       , fabric_data_to_bist_o12                                  => fabric_data_to_bist_o(11)
       , fabric_data_to_bist_o13                                  => fabric_data_to_bist_o(12)
       , fabric_data_to_bist_o14                                  => fabric_data_to_bist_o(13)
       , fabric_data_to_bist_o15                                  => fabric_data_to_bist_o(14)
       , fabric_data_to_bist_o16                                  => fabric_data_to_bist_o(15)
       , fabric_data_to_bist_o17                                  => fabric_data_to_bist_o(16)
       , fabric_data_to_bist_o18                                  => fabric_data_to_bist_o(17)
       , fabric_data_to_bist_o19                                  => fabric_data_to_bist_o(18)
       , fabric_data_to_bist_o20                                  => fabric_data_to_bist_o(19)
       , fabric_data_to_bist_o21                                  => fabric_data_to_bist_o(20)
       , fabric_data_to_bist_o22                                  => fabric_data_to_bist_o(21)
       , fabric_data_to_bist_o23                                  => fabric_data_to_bist_o(22)
       , fabric_data_to_bist_o24                                  => fabric_data_to_bist_o(23)
       , fabric_otp_user_startword_o1                             => fabric_otp_user_startword_o(0)
       , fabric_otp_user_startword_o2                             => fabric_otp_user_startword_o(1)
       , fabric_otp_user_startword_o3                             => fabric_otp_user_startword_o(2)
       , fabric_otp_user_startword_o4                             => fabric_otp_user_startword_o(3)
       , fabric_otp_user_startword_o5                             => fabric_otp_user_startword_o(4)
       , fabric_otp_user_startword_o6                             => fabric_otp_user_startword_o(5)
       , fabric_otp_user_startword_o7                             => fabric_otp_user_startword_o(6)
       , fabric_otp_user_startword_o8                             => fabric_otp_user_startword_o(7)
       , fabric_otp_user_startword_o9                             => fabric_otp_user_startword_o(8)
       , fabric_otp_user_startword_o10                            => fabric_otp_user_startword_o(9)
       , fabric_otp_user_startword_o11                            => fabric_otp_user_startword_o(10)
       , fabric_otp_user_startword_o12                            => fabric_otp_user_startword_o(11)
       , fabric_otp_user_startword_o13                            => fabric_otp_user_startword_o(12)
       , fabric_otp_user_startword_o14                            => fabric_otp_user_startword_o(13)
       , fabric_otp_user_startword_o15                            => fabric_otp_user_startword_o(14)
       , fabric_otp_user_startword_o16                            => fabric_otp_user_startword_o(15)
       , fabric_ahb_direct_data_o1                                => fabric_ahb_direct_data_o(0)
       , fabric_ahb_direct_data_o2                                => fabric_ahb_direct_data_o(1)
       , fabric_ahb_direct_data_o3                                => fabric_ahb_direct_data_o(2)
       , fabric_ahb_direct_data_o4                                => fabric_ahb_direct_data_o(3)
       , fabric_ahb_direct_data_o5                                => fabric_ahb_direct_data_o(4)
       , fabric_ahb_direct_data_o6                                => fabric_ahb_direct_data_o(5)
       , fabric_ahb_direct_data_o7                                => fabric_ahb_direct_data_o(6)
       , fabric_ahb_direct_data_o8                                => fabric_ahb_direct_data_o(7)
       , fabric_ahb_direct_data_o9                                => fabric_ahb_direct_data_o(8)
       , fabric_ahb_direct_data_o10                               => fabric_ahb_direct_data_o(9)
       , fabric_ahb_direct_data_o11                               => fabric_ahb_direct_data_o(10)
       , fabric_ahb_direct_data_o12                               => fabric_ahb_direct_data_o(11)
       , fabric_ahb_direct_data_o13                               => fabric_ahb_direct_data_o(12)
       , fabric_ahb_direct_data_o14                               => fabric_ahb_direct_data_o(13)
       , fabric_ahb_direct_data_o15                               => fabric_ahb_direct_data_o(14)
       , fabric_ahb_direct_data_o16                               => fabric_ahb_direct_data_o(15)
       , fabric_ahb_direct_data_o17                               => fabric_ahb_direct_data_o(16)
       , fabric_ahb_direct_data_o18                               => fabric_ahb_direct_data_o(17)
       , fabric_ahb_direct_data_o19                               => fabric_ahb_direct_data_o(18)
       , fabric_ahb_direct_data_o20                               => fabric_ahb_direct_data_o(19)
       , fabric_ahb_direct_data_o21                               => fabric_ahb_direct_data_o(20)
       , fabric_ahb_direct_data_o22                               => fabric_ahb_direct_data_o(21)
       , fabric_ahb_direct_data_o23                               => fabric_ahb_direct_data_o(22)
       , fabric_ahb_direct_data_o24                               => fabric_ahb_direct_data_o(23)
       , fabric_ahb_direct_data_o25                               => fabric_ahb_direct_data_o(24)
       , fabric_ahb_direct_data_o26                               => fabric_ahb_direct_data_o(25)
       , fabric_ahb_direct_data_o27                               => fabric_ahb_direct_data_o(26)
       , fabric_ahb_direct_data_o28                               => fabric_ahb_direct_data_o(27)
       , fabric_ahb_direct_data_o29                               => fabric_ahb_direct_data_o(28)
       , fabric_ahb_direct_data_o30                               => fabric_ahb_direct_data_o(29)
       , fabric_ahb_direct_data_o31                               => fabric_ahb_direct_data_o(30)
       , fabric_ahb_direct_data_o32                               => fabric_ahb_direct_data_o(31)
       , fabric_parusr_data_o1                                    => fabric_parusr_data_o(0)
       , fabric_parusr_data_o2                                    => fabric_parusr_data_o(1)
       , fabric_parusr_data_o3                                    => fabric_parusr_data_o(2)
       , fabric_parusr_data_o4                                    => fabric_parusr_data_o(3)
       , fabric_parusr_data_o5                                    => fabric_parusr_data_o(4)
       , fabric_parusr_data_o6                                    => fabric_parusr_data_o(5)
       , fabric_parusr_data_o7                                    => fabric_parusr_data_o(6)
       , fabric_parusr_data_o8                                    => fabric_parusr_data_o(7)
       , fabric_parusr_data_o9                                    => fabric_parusr_data_o(8)
       , fabric_parusr_data_o10                                   => fabric_parusr_data_o(9)
       , fabric_parusr_data_o11                                   => fabric_parusr_data_o(10)
       , fabric_parusr_data_o12                                   => fabric_parusr_data_o(11)
       , fabric_parusr_data_o13                                   => fabric_parusr_data_o(12)
       , fabric_parusr_data_o14                                   => fabric_parusr_data_o(13)
       , fabric_parusr_data_o15                                   => fabric_parusr_data_o(14)
       , fabric_parusr_data_o16                                   => fabric_parusr_data_o(15)
       , fabric_debug_otp_reload_err_o                            => fabric_debug_otp_reload_err_o
       , fabric_cfg_fabric_user_unmask_o                          => fabric_cfg_fabric_user_unmask_o
       , fabric_decoder_init_ready_o                              => fabric_decoder_init_ready_o
       , fabric_global_chip_status_o1                             => fabric_global_chip_status_o(0)
       , fabric_global_chip_status_o2                             => fabric_global_chip_status_o(1)
       , fabric_global_chip_status_o3                             => fabric_global_chip_status_o(2)
       , fabric_debug_security_boot_done_o                        => fabric_debug_security_boot_done_o
       , fabric_otp_user_calibrated_o                             => fabric_otp_user_calibrated_o
       , fabric_fuse_status_o1                                    => fabric_fuse_status_o(0)
       , fabric_fuse_status_o2                                    => fabric_fuse_status_o(1)
       , fabric_fuse_status_o3                                    => fabric_fuse_status_o(2)
       , fabric_otp_apb_rdata_o1                                  => fabric_otp_apb_rdata_o(0)
       , fabric_otp_apb_rdata_o2                                  => fabric_otp_apb_rdata_o(1)
       , fabric_otp_apb_rdata_o3                                  => fabric_otp_apb_rdata_o(2)
       , fabric_otp_apb_rdata_o4                                  => fabric_otp_apb_rdata_o(3)
       , fabric_otp_apb_rdata_o5                                  => fabric_otp_apb_rdata_o(4)
       , fabric_otp_apb_rdata_o6                                  => fabric_otp_apb_rdata_o(5)
       , fabric_otp_apb_rdata_o7                                  => fabric_otp_apb_rdata_o(6)
       , fabric_otp_apb_rdata_o8                                  => fabric_otp_apb_rdata_o(7)
       , fabric_otp_apb_rdata_o9                                  => fabric_otp_apb_rdata_o(8)
       , fabric_otp_apb_rdata_o10                                 => fabric_otp_apb_rdata_o(9)
       , fabric_otp_apb_rdata_o11                                 => fabric_otp_apb_rdata_o(10)
       , fabric_otp_apb_rdata_o12                                 => fabric_otp_apb_rdata_o(11)
       , fabric_otp_apb_rdata_o13                                 => fabric_otp_apb_rdata_o(12)
       , fabric_otp_apb_rdata_o14                                 => fabric_otp_apb_rdata_o(13)
       , fabric_otp_apb_rdata_o15                                 => fabric_otp_apb_rdata_o(14)
       , fabric_otp_apb_rdata_o16                                 => fabric_otp_apb_rdata_o(15)
       , fabric_otp_apb_rdata_o17                                 => fabric_otp_apb_rdata_o(16)
       , fabric_otp_apb_rdata_o18                                 => fabric_otp_apb_rdata_o(17)
       , fabric_otp_apb_rdata_o19                                 => fabric_otp_apb_rdata_o(18)
       , fabric_otp_apb_rdata_o20                                 => fabric_otp_apb_rdata_o(19)
       , fabric_otp_apb_rdata_o21                                 => fabric_otp_apb_rdata_o(20)
       , fabric_otp_apb_rdata_o22                                 => fabric_otp_apb_rdata_o(21)
       , fabric_otp_apb_rdata_o23                                 => fabric_otp_apb_rdata_o(22)
       , fabric_otp_apb_rdata_o24                                 => fabric_otp_apb_rdata_o(23)
       , fabric_otp_apb_rdata_o25                                 => fabric_otp_apb_rdata_o(24)
       , fabric_otp_apb_rdata_o26                                 => fabric_otp_apb_rdata_o(25)
       , fabric_otp_apb_rdata_o27                                 => fabric_otp_apb_rdata_o(26)
       , fabric_otp_apb_rdata_o28                                 => fabric_otp_apb_rdata_o(27)
       , fabric_otp_apb_rdata_o29                                 => fabric_otp_apb_rdata_o(28)
       , fabric_otp_apb_rdata_o30                                 => fabric_otp_apb_rdata_o(29)
       , fabric_otp_apb_rdata_o31                                 => fabric_otp_apb_rdata_o(30)
       , fabric_otp_apb_rdata_o32                                 => fabric_otp_apb_rdata_o(31)
       , fabric_jtag_tms_o                                        => fabric_jtag_tms_o
       , fabric_debug_bsec_core_status_o1                         => fabric_debug_bsec_core_status_o(0)
       , fabric_debug_bsec_core_status_o2                         => fabric_debug_bsec_core_status_o(1)
       , fabric_debug_bsec_core_status_o3                         => fabric_debug_bsec_core_status_o(2)
       , fabric_debug_bsec_core_status_o4                         => fabric_debug_bsec_core_status_o(3)
       , fabric_debug_bsec_core_status_o5                         => fabric_debug_bsec_core_status_o(4)
       , fabric_debug_bsec_core_status_o6                         => fabric_debug_bsec_core_status_o(5)
       , fabric_debug_bsec_core_status_o7                         => fabric_debug_bsec_core_status_o(6)
       , fabric_debug_bsec_core_status_o8                         => fabric_debug_bsec_core_status_o(7)
       , fabric_debug_bsec_core_status_o9                         => fabric_debug_bsec_core_status_o(8)
       , fabric_debug_bsec_core_status_o10                        => fabric_debug_bsec_core_status_o(9)
       , fabric_debug_bsec_core_status_o11                        => fabric_debug_bsec_core_status_o(10)
       , fabric_debug_bsec_core_status_o12                        => fabric_debug_bsec_core_status_o(11)
       , fabric_debug_bsec_core_status_o13                        => fabric_debug_bsec_core_status_o(12)
       , fabric_debug_bsec_core_status_o14                        => fabric_debug_bsec_core_status_o(13)
       , fabric_debug_bsec_core_status_o15                        => fabric_debug_bsec_core_status_o(14)
       , fabric_debug_bsec_core_status_o16                        => fabric_debug_bsec_core_status_o(15)
       , fabric_debug_bsec_core_status_o17                        => fabric_debug_bsec_core_status_o(16)
       , fabric_debug_bsec_core_status_o18                        => fabric_debug_bsec_core_status_o(17)
       , fabric_debug_bsec_core_status_o19                        => fabric_debug_bsec_core_status_o(18)
       , fabric_debug_bsec_core_status_o20                        => fabric_debug_bsec_core_status_o(19)
       , fabric_debug_bsec_core_status_o21                        => fabric_debug_bsec_core_status_o(20)
       , fabric_debug_bsec_core_status_o22                        => fabric_debug_bsec_core_status_o(21)
       , fabric_debug_bsec_core_status_o23                        => fabric_debug_bsec_core_status_o(22)
       , fabric_debug_bsec_core_status_o24                        => fabric_debug_bsec_core_status_o(23)
       , fabric_debug_bsec_core_status_o25                        => fabric_debug_bsec_core_status_o(24)
       , fabric_debug_bsec_core_status_o26                        => fabric_debug_bsec_core_status_o(25)
       , fabric_debug_bsec_core_status_o27                        => fabric_debug_bsec_core_status_o(26)
       , fabric_debug_bsec_core_status_o28                        => fabric_debug_bsec_core_status_o(27)
       , fabric_debug_bsec_core_status_o29                        => fabric_debug_bsec_core_status_o(28)
       , fabric_debug_bsec_core_status_o30                        => fabric_debug_bsec_core_status_o(29)
       , fabric_debug_bsec_core_status_o31                        => fabric_debug_bsec_core_status_o(30)
       , fabric_debug_bsec_core_status_o32                        => fabric_debug_bsec_core_status_o(31)
       , fabric_mrepair_fuse_bist1fail_o1                         => fabric_mrepair_fuse_bist1fail_o(0)
       , fabric_mrepair_fuse_bist1fail_o2                         => fabric_mrepair_fuse_bist1fail_o(1)
       , fabric_mrepair_fuse_bist1fail_o3                         => fabric_mrepair_fuse_bist1fail_o(2)
       , fabric_mrepair_fuse_bist1fail_o4                         => fabric_mrepair_fuse_bist1fail_o(3)
       , fabric_mrepair_fuse_bist1fail_o5                         => fabric_mrepair_fuse_bist1fail_o(4)
       , fabric_mrepair_fuse_bist1fail_o6                         => fabric_mrepair_fuse_bist1fail_o(5)
       , fabric_mrepair_fuse_bist1fail_o7                         => fabric_mrepair_fuse_bist1fail_o(6)
       , fabric_mrepair_fuse_bist1fail_o8                         => fabric_mrepair_fuse_bist1fail_o(7)
       , fabric_flag_ready_o                                      => fabric_flag_ready_o
       , fabric_mrepair_fuse_dout_o1                              => fabric_mrepair_fuse_dout_o(0)
       , fabric_mrepair_fuse_dout_o2                              => fabric_mrepair_fuse_dout_o(1)
       , fabric_mrepair_fuse_dout_o3                              => fabric_mrepair_fuse_dout_o(2)
       , fabric_mrepair_fuse_dout_o4                              => fabric_mrepair_fuse_dout_o(3)
       , fabric_mrepair_fuse_dout_o5                              => fabric_mrepair_fuse_dout_o(4)
       , fabric_mrepair_fuse_dout_o6                              => fabric_mrepair_fuse_dout_o(5)
       , fabric_mrepair_fuse_dout_o7                              => fabric_mrepair_fuse_dout_o(6)
       , fabric_mrepair_fuse_dout_o8                              => fabric_mrepair_fuse_dout_o(7)
       , fabric_mrepair_fuse_dout_o9                              => fabric_mrepair_fuse_dout_o(8)
       , fabric_mrepair_fuse_dout_o10                             => fabric_mrepair_fuse_dout_o(9)
       , fabric_mrepair_fuse_dout_o11                             => fabric_mrepair_fuse_dout_o(10)
       , fabric_mrepair_fuse_dout_o12                             => fabric_mrepair_fuse_dout_o(11)
       , fabric_mrepair_fuse_dout_o13                             => fabric_mrepair_fuse_dout_o(12)
       , fabric_mrepair_fuse_dout_o14                             => fabric_mrepair_fuse_dout_o(13)
       , fabric_mrepair_fuse_dout_o15                             => fabric_mrepair_fuse_dout_o(14)
       , fabric_mrepair_fuse_dout_o16                             => fabric_mrepair_fuse_dout_o(15)
       , fabric_mrepair_fuse_dout_o17                             => fabric_mrepair_fuse_dout_o(16)
       , fabric_mrepair_fuse_dout_o18                             => fabric_mrepair_fuse_dout_o(17)
       , fabric_mrepair_fuse_dout_o19                             => fabric_mrepair_fuse_dout_o(18)
       , fabric_mrepair_fuse_dout_o20                             => fabric_mrepair_fuse_dout_o(19)
       , fabric_mrepair_fuse_dout_o21                             => fabric_mrepair_fuse_dout_o(20)
       , fabric_mrepair_fuse_dout_o22                             => fabric_mrepair_fuse_dout_o(21)
       , fabric_mrepair_fuse_dout_o23                             => fabric_mrepair_fuse_dout_o(22)
       , fabric_mrepair_fuse_dout_o24                             => fabric_mrepair_fuse_dout_o(23)
       , fabric_mrepair_fuse_dout_o25                             => fabric_mrepair_fuse_dout_o(24)
       , fabric_mrepair_fuse_dout_o26                             => fabric_mrepair_fuse_dout_o(25)
       , fabric_mrepair_fuse_dout_o27                             => fabric_mrepair_fuse_dout_o(26)
       , fabric_mrepair_fuse_dout_o28                             => fabric_mrepair_fuse_dout_o(27)
       , fabric_mrepair_fuse_dout_o29                             => fabric_mrepair_fuse_dout_o(28)
       , fabric_mrepair_fuse_dout_o30                             => fabric_mrepair_fuse_dout_o(29)
       , fabric_mrepair_fuse_dout_o31                             => fabric_mrepair_fuse_dout_o(30)
       , fabric_mrepair_fuse_dout_o32                             => fabric_mrepair_fuse_dout_o(31)
       , fabric_mrepair_fuse_dout_o33                             => fabric_mrepair_fuse_dout_o(32)
       , fabric_mrepair_fuse_dout_o34                             => fabric_mrepair_fuse_dout_o(33)
       , fabric_mrepair_fuse_dout_o35                             => fabric_mrepair_fuse_dout_o(34)
       , fabric_mrepair_fuse_dout_o36                             => fabric_mrepair_fuse_dout_o(35)
       , fabric_mrepair_fuse_dout_o37                             => fabric_mrepair_fuse_dout_o(36)
       , fabric_mrepair_fuse_dout_o38                             => fabric_mrepair_fuse_dout_o(37)
       , fabric_mrepair_fuse_dout_o39                             => fabric_mrepair_fuse_dout_o(38)
       , fabric_mrepair_fuse_dout_o40                             => fabric_mrepair_fuse_dout_o(39)
       , fabric_mrepair_fuse_dout_o41                             => fabric_mrepair_fuse_dout_o(40)
       , fabric_debug_rst_soft_o                                  => fabric_debug_rst_soft_o
       , fabric_otp_user_ack_o                                    => fabric_otp_user_ack_o
       , fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o  => fabric_mrepair_fuse_prg_block_space_read_error_flag_q_o
       , fabric_shift_en_to_bist_o1                               => fabric_shift_en_to_bist_o(0)
       , fabric_shift_en_to_bist_o2                               => fabric_shift_en_to_bist_o(1)
       , fabric_shift_en_to_bist_o3                               => fabric_shift_en_to_bist_o(2)
       , fabric_shift_en_to_bist_o4                               => fabric_shift_en_to_bist_o(3)
       , fabric_shift_en_to_bist_o5                               => fabric_shift_en_to_bist_o(4)
       , fabric_shift_en_to_bist_o6                               => fabric_shift_en_to_bist_o(5)
       , fabric_shift_en_to_bist_o7                               => fabric_shift_en_to_bist_o(6)
       , fabric_shift_en_to_bist_o8                               => fabric_shift_en_to_bist_o(7)
       , fabric_shift_en_to_bist_o9                               => fabric_shift_en_to_bist_o(8)
       , fabric_shift_en_to_bist_o10                              => fabric_shift_en_to_bist_o(9)
       , fabric_shift_en_to_bist_o11                              => fabric_shift_en_to_bist_o(10)
       , fabric_shift_en_to_bist_o12                              => fabric_shift_en_to_bist_o(11)
       , fabric_shift_en_to_bist_o13                              => fabric_shift_en_to_bist_o(12)
       , fabric_shift_en_to_bist_o14                              => fabric_shift_en_to_bist_o(13)
       , fabric_shift_en_to_bist_o15                              => fabric_shift_en_to_bist_o(14)
       , fabric_shift_en_to_bist_o16                              => fabric_shift_en_to_bist_o(15)
       , fabric_shift_en_to_bist_o17                              => fabric_shift_en_to_bist_o(16)
       , fabric_shift_en_to_bist_o18                              => fabric_shift_en_to_bist_o(17)
       , fabric_shift_en_to_bist_o19                              => fabric_shift_en_to_bist_o(18)
       , fabric_shift_en_to_bist_o20                              => fabric_shift_en_to_bist_o(19)
       , fabric_shift_en_to_bist_o21                              => fabric_shift_en_to_bist_o(20)
       , fabric_shift_en_to_bist_o22                              => fabric_shift_en_to_bist_o(21)
       , fabric_shift_en_to_bist_o23                              => fabric_shift_en_to_bist_o(22)
       , fabric_shift_en_to_bist_o24                              => fabric_shift_en_to_bist_o(23)
       , fabric_sif_reg_en_to_bist_o1                             => fabric_sif_reg_en_to_bist_o(0)
       , fabric_sif_reg_en_to_bist_o2                             => fabric_sif_reg_en_to_bist_o(1)
       , fabric_sif_reg_en_to_bist_o3                             => fabric_sif_reg_en_to_bist_o(2)
       , fabric_sif_reg_en_to_bist_o4                             => fabric_sif_reg_en_to_bist_o(3)
       , fabric_sif_reg_en_to_bist_o5                             => fabric_sif_reg_en_to_bist_o(4)
       , fabric_sif_reg_en_to_bist_o6                             => fabric_sif_reg_en_to_bist_o(5)
       , fabric_sif_reg_en_to_bist_o7                             => fabric_sif_reg_en_to_bist_o(6)
       , fabric_sif_reg_en_to_bist_o8                             => fabric_sif_reg_en_to_bist_o(7)
       , fabric_sif_reg_en_to_bist_o9                             => fabric_sif_reg_en_to_bist_o(8)
       , fabric_sif_reg_en_to_bist_o10                            => fabric_sif_reg_en_to_bist_o(9)
       , fabric_sif_reg_en_to_bist_o11                            => fabric_sif_reg_en_to_bist_o(10)
       , fabric_sif_reg_en_to_bist_o12                            => fabric_sif_reg_en_to_bist_o(11)
       , fabric_sif_reg_en_to_bist_o13                            => fabric_sif_reg_en_to_bist_o(12)
       , fabric_sif_reg_en_to_bist_o14                            => fabric_sif_reg_en_to_bist_o(13)
       , fabric_sif_reg_en_to_bist_o15                            => fabric_sif_reg_en_to_bist_o(14)
       , fabric_sif_reg_en_to_bist_o16                            => fabric_sif_reg_en_to_bist_o(15)
       , fabric_sif_reg_en_to_bist_o17                            => fabric_sif_reg_en_to_bist_o(16)
       , fabric_sif_reg_en_to_bist_o18                            => fabric_sif_reg_en_to_bist_o(17)
       , fabric_sif_reg_en_to_bist_o19                            => fabric_sif_reg_en_to_bist_o(18)
       , fabric_sif_reg_en_to_bist_o20                            => fabric_sif_reg_en_to_bist_o(19)
       , fabric_sif_reg_en_to_bist_o21                            => fabric_sif_reg_en_to_bist_o(20)
       , fabric_sif_reg_en_to_bist_o22                            => fabric_sif_reg_en_to_bist_o(21)
       , fabric_sif_reg_en_to_bist_o23                            => fabric_sif_reg_en_to_bist_o(22)
       , fabric_sif_reg_en_to_bist_o24                            => fabric_sif_reg_en_to_bist_o(23)
       , fabric_sif_reg_en_to_bist_o25                            => fabric_sif_reg_en_to_bist_o(24)
       , fabric_sif_reg_en_to_bist_o26                            => fabric_sif_reg_en_to_bist_o(25)
       , fabric_sif_reg_en_to_bist_o27                            => fabric_sif_reg_en_to_bist_o(26)
       , fabric_sif_reg_en_to_bist_o28                            => fabric_sif_reg_en_to_bist_o(27)
       , fabric_sif_reg_en_to_bist_o29                            => fabric_sif_reg_en_to_bist_o(28)
       , fabric_sif_reg_en_to_bist_o30                            => fabric_sif_reg_en_to_bist_o(29)
       , fabric_sif_reg_en_to_bist_o31                            => fabric_sif_reg_en_to_bist_o(30)
       , fabric_sif_reg_en_to_bist_o32                            => fabric_sif_reg_en_to_bist_o(31)
       , fabric_sif_reg_en_to_bist_o33                            => fabric_sif_reg_en_to_bist_o(32)
       , fabric_sif_reg_en_to_bist_o34                            => fabric_sif_reg_en_to_bist_o(33)
       , fabric_sif_reg_en_to_bist_o35                            => fabric_sif_reg_en_to_bist_o(34)
       , fabric_sif_reg_en_to_bist_o36                            => fabric_sif_reg_en_to_bist_o(35)
       , fabric_sif_reg_en_to_bist_o37                            => fabric_sif_reg_en_to_bist_o(36)
       , fabric_sif_reg_en_to_bist_o38                            => fabric_sif_reg_en_to_bist_o(37)
       , fabric_sif_reg_en_to_bist_o39                            => fabric_sif_reg_en_to_bist_o(38)
       , fabric_sif_reg_en_to_bist_o40                            => fabric_sif_reg_en_to_bist_o(39)
       , fabric_sif_reg_en_to_bist_o41                            => fabric_sif_reg_en_to_bist_o(40)
       , fabric_sif_reg_en_to_bist_o42                            => fabric_sif_reg_en_to_bist_o(41)
       , fabric_sif_reg_en_to_bist_o43                            => fabric_sif_reg_en_to_bist_o(42)
       , fabric_sif_reg_en_to_bist_o44                            => fabric_sif_reg_en_to_bist_o(43)
       , fabric_sif_reg_en_to_bist_o45                            => fabric_sif_reg_en_to_bist_o(44)
       , fabric_sif_reg_en_to_bist_o46                            => fabric_sif_reg_en_to_bist_o(45)
       , fabric_sif_reg_en_to_bist_o47                            => fabric_sif_reg_en_to_bist_o(46)
       , fabric_sif_reg_en_to_bist_o48                            => fabric_sif_reg_en_to_bist_o(47)
       , fabric_sif_reg_en_to_bist_o49                            => fabric_sif_reg_en_to_bist_o(48)
       , fabric_sif_reg_en_to_bist_o50                            => fabric_sif_reg_en_to_bist_o(49)
       , fabric_sif_reg_en_to_bist_o51                            => fabric_sif_reg_en_to_bist_o(50)
       , fabric_sif_reg_en_to_bist_o52                            => fabric_sif_reg_en_to_bist_o(51)
       , fabric_sif_reg_en_to_bist_o53                            => fabric_sif_reg_en_to_bist_o(52)
       , fabric_sif_reg_en_to_bist_o54                            => fabric_sif_reg_en_to_bist_o(53)
       , fabric_sif_reg_en_to_bist_o55                            => fabric_sif_reg_en_to_bist_o(54)
       , fabric_sif_reg_en_to_bist_o56                            => fabric_sif_reg_en_to_bist_o(55)
       , fabric_sif_reg_en_to_bist_o57                            => fabric_sif_reg_en_to_bist_o(56)
       , fabric_sif_reg_en_to_bist_o58                            => fabric_sif_reg_en_to_bist_o(57)
       , fabric_sif_reg_en_to_bist_o59                            => fabric_sif_reg_en_to_bist_o(58)
       , fabric_sif_reg_en_to_bist_o60                            => fabric_sif_reg_en_to_bist_o(59)
       , fabric_sif_reg_en_to_bist_o61                            => fabric_sif_reg_en_to_bist_o(60)
       , fabric_sif_reg_en_to_bist_o62                            => fabric_sif_reg_en_to_bist_o(61)
       , fabric_sif_reg_en_to_bist_o63                            => fabric_sif_reg_en_to_bist_o(62)
       , fabric_sif_reg_en_to_bist_o64                            => fabric_sif_reg_en_to_bist_o(63)
       , fabric_sif_reg_en_to_bist_o65                            => fabric_sif_reg_en_to_bist_o(64)
       , fabric_sif_reg_en_to_bist_o66                            => fabric_sif_reg_en_to_bist_o(65)
       , fabric_sif_reg_en_to_bist_o67                            => fabric_sif_reg_en_to_bist_o(66)
       , fabric_sif_reg_en_to_bist_o68                            => fabric_sif_reg_en_to_bist_o(67)
       , fabric_sif_reg_en_to_bist_o69                            => fabric_sif_reg_en_to_bist_o(68)
       , fabric_sif_reg_en_to_bist_o70                            => fabric_sif_reg_en_to_bist_o(69)
       , fabric_sif_reg_en_to_bist_o71                            => fabric_sif_reg_en_to_bist_o(70)
       , fabric_sif_reg_en_to_bist_o72                            => fabric_sif_reg_en_to_bist_o(71)
       , fabric_sif_reg_en_to_bist_o73                            => fabric_sif_reg_en_to_bist_o(72)
       , fabric_sif_reg_en_to_bist_o74                            => fabric_sif_reg_en_to_bist_o(73)
       , fabric_sif_reg_en_to_bist_o75                            => fabric_sif_reg_en_to_bist_o(74)
       , fabric_sif_reg_en_to_bist_o76                            => fabric_sif_reg_en_to_bist_o(75)
       , fabric_sif_reg_en_to_bist_o77                            => fabric_sif_reg_en_to_bist_o(76)
       , fabric_sif_reg_en_to_bist_o78                            => fabric_sif_reg_en_to_bist_o(77)
       , fabric_sif_reg_en_to_bist_o79                            => fabric_sif_reg_en_to_bist_o(78)
       , fabric_sif_reg_en_to_bist_o80                            => fabric_sif_reg_en_to_bist_o(79)
       , fabric_sif_reg_en_to_bist_o81                            => fabric_sif_reg_en_to_bist_o(80)
       , fabric_sif_reg_en_to_bist_o82                            => fabric_sif_reg_en_to_bist_o(81)
       , fabric_sif_reg_en_to_bist_o83                            => fabric_sif_reg_en_to_bist_o(82)
       , fabric_sif_reg_en_to_bist_o84                            => fabric_sif_reg_en_to_bist_o(83)
       , fabric_sif_reg_en_to_bist_o85                            => fabric_sif_reg_en_to_bist_o(84)
       , fabric_sif_reg_en_to_bist_o86                            => fabric_sif_reg_en_to_bist_o(85)
       , fabric_sif_reg_en_to_bist_o87                            => fabric_sif_reg_en_to_bist_o(86)
       , fabric_sif_reg_en_to_bist_o88                            => fabric_sif_reg_en_to_bist_o(87)
       , fabric_sif_reg_en_to_bist_o89                            => fabric_sif_reg_en_to_bist_o(88)
       , fabric_sif_reg_en_to_bist_o90                            => fabric_sif_reg_en_to_bist_o(89)
       , fabric_sif_reg_en_to_bist_o91                            => fabric_sif_reg_en_to_bist_o(90)
       , fabric_sif_reg_en_to_bist_o92                            => fabric_sif_reg_en_to_bist_o(91)
       , fabric_sif_reg_en_to_bist_o93                            => fabric_sif_reg_en_to_bist_o(92)
       , fabric_sif_reg_en_to_bist_o94                            => fabric_sif_reg_en_to_bist_o(93)
       , fabric_sif_reg_en_to_bist_o95                            => fabric_sif_reg_en_to_bist_o(94)
       , fabric_sif_reg_en_to_bist_o96                            => fabric_sif_reg_en_to_bist_o(95)
       , fabric_sif_reg_en_to_bist_o97                            => fabric_sif_reg_en_to_bist_o(96)
       , fabric_sif_reg_en_to_bist_o98                            => fabric_sif_reg_en_to_bist_o(97)
       , fabric_sif_reg_en_to_bist_o99                            => fabric_sif_reg_en_to_bist_o(98)
       , fabric_sif_reg_en_to_bist_o100                           => fabric_sif_reg_en_to_bist_o(99)
       , fabric_sif_reg_en_to_bist_o101                           => fabric_sif_reg_en_to_bist_o(100)
       , fabric_sif_reg_en_to_bist_o102                           => fabric_sif_reg_en_to_bist_o(101)
       , fabric_sif_reg_en_to_bist_o103                           => fabric_sif_reg_en_to_bist_o(102)
       , fabric_sif_reg_en_to_bist_o104                           => fabric_sif_reg_en_to_bist_o(103)
       , fabric_sif_reg_en_to_bist_o105                           => fabric_sif_reg_en_to_bist_o(104)
       , fabric_sif_reg_en_to_bist_o106                           => fabric_sif_reg_en_to_bist_o(105)
       , fabric_sif_reg_en_to_bist_o107                           => fabric_sif_reg_en_to_bist_o(106)
       , fabric_sif_reg_en_to_bist_o108                           => fabric_sif_reg_en_to_bist_o(107)
       , fabric_sif_reg_en_to_bist_o109                           => fabric_sif_reg_en_to_bist_o(108)
       , fabric_sif_reg_en_to_bist_o110                           => fabric_sif_reg_en_to_bist_o(109)
       , fabric_sif_reg_en_to_bist_o111                           => fabric_sif_reg_en_to_bist_o(110)
       , fabric_sif_reg_en_to_bist_o112                           => fabric_sif_reg_en_to_bist_o(111)
       , fabric_sif_reg_en_to_bist_o113                           => fabric_sif_reg_en_to_bist_o(112)
       , fabric_sif_reg_en_to_bist_o114                           => fabric_sif_reg_en_to_bist_o(113)
       , fabric_sif_reg_en_to_bist_o115                           => fabric_sif_reg_en_to_bist_o(114)
       , fabric_sif_reg_en_to_bist_o116                           => fabric_sif_reg_en_to_bist_o(115)
       , fabric_sif_reg_en_to_bist_o117                           => fabric_sif_reg_en_to_bist_o(116)
       , fabric_sif_reg_en_to_bist_o118                           => fabric_sif_reg_en_to_bist_o(117)
       , fabric_sif_reg_en_to_bist_o119                           => fabric_sif_reg_en_to_bist_o(118)
       , fabric_sif_reg_en_to_bist_o120                           => fabric_sif_reg_en_to_bist_o(119)
       , fabric_debug_otp_manager_read_otp_o                      => fabric_debug_otp_manager_read_otp_o
       , fabric_otp_user_sec_o                                    => fabric_otp_user_sec_o
       , fabric_otp_user_wlromout_o1                              => fabric_otp_user_wlromout_o(0)
       , fabric_otp_user_wlromout_o2                              => fabric_otp_user_wlromout_o(1)
       , fabric_otp_user_wlromout_o3                              => fabric_otp_user_wlromout_o(2)
       , fabric_otp_user_wlromout_o4                              => fabric_otp_user_wlromout_o(3)
       , fabric_otp_user_wlromout_o5                              => fabric_otp_user_wlromout_o(4)
       , fabric_otp_user_wlromout_o6                              => fabric_otp_user_wlromout_o(5)
       , fabric_otp_user_wlromout_o7                              => fabric_otp_user_wlromout_o(6)
       , fabric_otp_user_wlromout_o8                              => fabric_otp_user_wlromout_o(7)
       , fabric_otp_user_wlromout_o9                              => fabric_otp_user_wlromout_o(8)
       , fabric_otp_user_wlromout_o10                             => fabric_otp_user_wlromout_o(9)
       , fabric_mrepair_fuse_bend1_o                              => fabric_mrepair_fuse_bend1_o
       , fabric_mrepair_fuse_flagstate_o1                         => fabric_mrepair_fuse_flagstate_o(0)
       , fabric_mrepair_fuse_flagstate_o2                         => fabric_mrepair_fuse_flagstate_o(1)
       , fabric_mrepair_fuse_flagstate_o3                         => fabric_mrepair_fuse_flagstate_o(2)
       , fabric_mrepair_fuse_flagstate_o4                         => fabric_mrepair_fuse_flagstate_o(3)
       , fabric_system_data_from_mem_bist_o1                      => fabric_system_data_from_mem_bist_o(0)
       , fabric_system_data_from_mem_bist_o2                      => fabric_system_data_from_mem_bist_o(1)
       , fabric_system_data_from_mem_bist_o3                      => fabric_system_data_from_mem_bist_o(2)
       , fabric_system_data_from_mem_bist_o4                      => fabric_system_data_from_mem_bist_o(3)
       , fabric_system_data_from_mem_bist_o5                      => fabric_system_data_from_mem_bist_o(4)
       , fabric_system_data_from_mem_bist_o6                      => fabric_system_data_from_mem_bist_o(5)
       , fabric_system_data_from_mem_bist_o7                      => fabric_system_data_from_mem_bist_o(6)
       , fabric_system_data_from_mem_bist_o8                      => fabric_system_data_from_mem_bist_o(7)
       , fabric_system_data_from_mem_bist_o9                      => fabric_system_data_from_mem_bist_o(8)
       , fabric_system_data_from_mem_bist_o10                     => fabric_system_data_from_mem_bist_o(9)
       , fabric_system_data_from_mem_bist_o11                     => fabric_system_data_from_mem_bist_o(10)
       , fabric_system_data_from_mem_bist_o12                     => fabric_system_data_from_mem_bist_o(11)
       , fabric_system_data_from_mem_bist_o13                     => fabric_system_data_from_mem_bist_o(12)
       , fabric_system_data_from_mem_bist_o14                     => fabric_system_data_from_mem_bist_o(13)
       , fabric_system_data_from_mem_bist_o15                     => fabric_system_data_from_mem_bist_o(14)
       , fabric_system_data_from_mem_bist_o16                     => fabric_system_data_from_mem_bist_o(15)
       , fabric_system_data_from_mem_bist_o17                     => fabric_system_data_from_mem_bist_o(16)
       , fabric_system_data_from_mem_bist_o18                     => fabric_system_data_from_mem_bist_o(17)
       , fabric_system_data_from_mem_bist_o19                     => fabric_system_data_from_mem_bist_o(18)
       , fabric_system_data_from_mem_bist_o20                     => fabric_system_data_from_mem_bist_o(19)
       , fabric_system_data_from_mem_bist_o21                     => fabric_system_data_from_mem_bist_o(20)
       , fabric_system_data_from_mem_bist_o22                     => fabric_system_data_from_mem_bist_o(21)
       , fabric_system_data_from_mem_bist_o23                     => fabric_system_data_from_mem_bist_o(22)
       , fabric_system_data_from_mem_bist_o24                     => fabric_system_data_from_mem_bist_o(23)
       , fabric_direct_data_o1                                    => fabric_direct_data_o(0)
       , fabric_direct_data_o2                                    => fabric_direct_data_o(1)
       , fabric_direct_data_o3                                    => fabric_direct_data_o(2)
       , fabric_direct_data_o4                                    => fabric_direct_data_o(3)
       , fabric_direct_data_o5                                    => fabric_direct_data_o(4)
       , fabric_direct_data_o6                                    => fabric_direct_data_o(5)
       , fabric_direct_data_o7                                    => fabric_direct_data_o(6)
       , fabric_direct_data_o8                                    => fabric_direct_data_o(7)
       , fabric_direct_data_o9                                    => fabric_direct_data_o(8)
       , fabric_direct_data_o10                                   => fabric_direct_data_o(9)
       , fabric_direct_data_o11                                   => fabric_direct_data_o(10)
       , fabric_direct_data_o12                                   => fabric_direct_data_o(11)
       , fabric_direct_data_o13                                   => fabric_direct_data_o(12)
       , fabric_direct_data_o14                                   => fabric_direct_data_o(13)
       , fabric_direct_data_o15                                   => fabric_direct_data_o(14)
       , fabric_direct_data_o16                                   => fabric_direct_data_o(15)
       , fabric_direct_data_o17                                   => fabric_direct_data_o(16)
       , fabric_direct_data_o18                                   => fabric_direct_data_o(17)
       , fabric_direct_data_o19                                   => fabric_direct_data_o(18)
       , fabric_direct_data_o20                                   => fabric_direct_data_o(19)
       , fabric_direct_data_o21                                   => fabric_direct_data_o(20)
       , fabric_direct_data_o22                                   => fabric_direct_data_o(21)
       , fabric_direct_data_o23                                   => fabric_direct_data_o(22)
       , fabric_direct_data_o24                                   => fabric_direct_data_o(23)
       , fabric_direct_data_o25                                   => fabric_direct_data_o(24)
       , fabric_direct_data_o26                                   => fabric_direct_data_o(25)
       , fabric_direct_data_o27                                   => fabric_direct_data_o(26)
       , fabric_direct_data_o28                                   => fabric_direct_data_o(27)
       , fabric_direct_data_o29                                   => fabric_direct_data_o(28)
       , fabric_direct_data_o30                                   => fabric_direct_data_o(29)
       , fabric_direct_data_o31                                   => fabric_direct_data_o(30)
       , fabric_direct_data_o32                                   => fabric_direct_data_o(31)
       , fabric_otp_user_bbad_o                                   => fabric_otp_user_bbad_o
       , fabric_user_read_cycle_o                                 => fabric_user_read_cycle_o
       , fabric_chip_status_o1                                    => fabric_chip_status_o(0)
       , fabric_chip_status_o2                                    => fabric_chip_status_o(1)
       , fabric_chip_status_o3                                    => fabric_chip_status_o(2)
       , fabric_chip_status_o4                                    => fabric_chip_status_o(3)
       , fabric_chip_status_o5                                    => fabric_chip_status_o(4)
       , fabric_chip_status_o6                                    => fabric_chip_status_o(5)
       , fabric_chip_status_o7                                    => fabric_chip_status_o(6)
       , fabric_chip_status_o8                                    => fabric_chip_status_o(7)
       , fabric_chip_status_o9                                    => fabric_chip_status_o(8)
       , fabric_chip_status_o10                                   => fabric_chip_status_o(9)
       , fabric_chip_status_o11                                   => fabric_chip_status_o(10)
       , fabric_chip_status_o12                                   => fabric_chip_status_o(11)
       , fabric_chip_status_o13                                   => fabric_chip_status_o(12)
       , fabric_chip_status_o14                                   => fabric_chip_status_o(13)
       , fabric_chip_status_o15                                   => fabric_chip_status_o(14)
       , fabric_chip_status_o16                                   => fabric_chip_status_o(15)
       , fabric_chip_status_o17                                   => fabric_chip_status_o(16)
       , fabric_chip_status_o18                                   => fabric_chip_status_o(17)
       , fabric_chip_status_o19                                   => fabric_chip_status_o(18)
       , fabric_chip_status_o20                                   => fabric_chip_status_o(19)
       , fabric_chip_status_o21                                   => fabric_chip_status_o(20)
       , fabric_chip_status_o22                                   => fabric_chip_status_o(21)
       , fabric_chip_status_o23                                   => fabric_chip_status_o(22)
       , fabric_chip_status_o24                                   => fabric_chip_status_o(23)
       , fabric_chip_status_o25                                   => fabric_chip_status_o(24)
       , fabric_chip_status_o26                                   => fabric_chip_status_o(25)
       , fabric_chip_status_o27                                   => fabric_chip_status_o(26)
       , fabric_chip_status_o28                                   => fabric_chip_status_o(27)
       , fabric_chip_status_o29                                   => fabric_chip_status_o(28)
       , fabric_chip_status_o30                                   => fabric_chip_status_o(29)
       , fabric_chip_status_o31                                   => fabric_chip_status_o(30)
       , fabric_chip_status_o32                                   => fabric_chip_status_o(31)
       , fabric_chip_status_o33                                   => fabric_chip_status_o(32)
       , fabric_chip_status_o34                                   => fabric_chip_status_o(33)
       , fabric_chip_status_o35                                   => fabric_chip_status_o(34)
       , fabric_chip_status_o36                                   => fabric_chip_status_o(35)
       , fabric_chip_status_o37                                   => fabric_chip_status_o(36)
       , fabric_chip_status_o38                                   => fabric_chip_status_o(37)
       , fabric_chip_status_o39                                   => fabric_chip_status_o(38)
       , fabric_chip_status_o40                                   => fabric_chip_status_o(39)
       , fabric_chip_status_o41                                   => fabric_chip_status_o(40)
       , fabric_chip_status_o42                                   => fabric_chip_status_o(41)
       , fabric_chip_status_o43                                   => fabric_chip_status_o(42)
       , fabric_chip_status_o44                                   => fabric_chip_status_o(43)
       , fabric_chip_status_o45                                   => fabric_chip_status_o(44)
       , fabric_chip_status_o46                                   => fabric_chip_status_o(45)
       , fabric_chip_status_o47                                   => fabric_chip_status_o(46)
       , fabric_chip_status_o48                                   => fabric_chip_status_o(47)
       , fabric_chip_status_o49                                   => fabric_chip_status_o(48)
       , fabric_chip_status_o50                                   => fabric_chip_status_o(49)
       , fabric_chip_status_o51                                   => fabric_chip_status_o(50)
       , fabric_chip_status_o52                                   => fabric_chip_status_o(51)
       , fabric_chip_status_o53                                   => fabric_chip_status_o(52)
       , fabric_chip_status_o54                                   => fabric_chip_status_o(53)
       , fabric_chip_status_o55                                   => fabric_chip_status_o(54)
       , fabric_chip_status_o56                                   => fabric_chip_status_o(55)
       , fabric_chip_status_o57                                   => fabric_chip_status_o(56)
       , fabric_chip_status_o58                                   => fabric_chip_status_o(57)
       , fabric_chip_status_o59                                   => fabric_chip_status_o(58)
       , fabric_chip_status_o60                                   => fabric_chip_status_o(59)
       , fabric_chip_status_o61                                   => fabric_chip_status_o(60)
       , fabric_chip_status_o62                                   => fabric_chip_status_o(61)
       , fabric_chip_status_o63                                   => fabric_chip_status_o(62)
       , fabric_chip_status_o64                                   => fabric_chip_status_o(63)
       , fabric_chip_status_o65                                   => fabric_chip_status_o(64)
       , fabric_chip_status_o66                                   => fabric_chip_status_o(65)
       , fabric_chip_status_o67                                   => fabric_chip_status_o(66)
       , fabric_chip_status_o68                                   => fabric_chip_status_o(67)
       , fabric_chip_status_o69                                   => fabric_chip_status_o(68)
       , fabric_chip_status_o70                                   => fabric_chip_status_o(69)
       , fabric_chip_status_o71                                   => fabric_chip_status_o(70)
       , fabric_chip_status_o72                                   => fabric_chip_status_o(71)
       , fabric_mrepair_fuse_disturbed_o                          => fabric_mrepair_fuse_disturbed_o
       , fabric_debug_otpboot_state_o1                            => fabric_debug_otpboot_state_o(0)
       , fabric_debug_otpboot_state_o2                            => fabric_debug_otpboot_state_o(1)
       , fabric_debug_otpboot_state_o3                            => fabric_debug_otpboot_state_o(2)
       , fabric_pd_ready_o1                                       => fabric_pd_ready_o(0)
       , fabric_pd_ready_o2                                       => fabric_pd_ready_o(1)
       , fabric_pd_ready_o3                                       => fabric_pd_ready_o(2)
       , fabric_pd_ready_o4                                       => fabric_pd_ready_o(3)
       , fabric_pd_ready_o5                                       => fabric_pd_ready_o(4)
       , fabric_pd_ready_o6                                       => fabric_pd_ready_o(5)
       , fabric_pd_ready_o7                                       => fabric_pd_ready_o(6)
       , fabric_pd_ready_o8                                       => fabric_pd_ready_o(7)
       , fabric_pd_ready_o9                                       => fabric_pd_ready_o(8)
       , fabric_pd_ready_o10                                      => fabric_pd_ready_o(9)
       , fabric_pd_ready_o11                                      => fabric_pd_ready_o(10)
       , fabric_pd_ready_o12                                      => fabric_pd_ready_o(11)
       , fabric_pd_ready_o13                                      => fabric_pd_ready_o(12)
       , fabric_pd_ready_o14                                      => fabric_pd_ready_o(13)
       , fabric_pd_ready_o15                                      => fabric_pd_ready_o(14)
       , fabric_pd_ready_o16                                      => fabric_pd_ready_o(15)
       , fabric_pd_ready_o17                                      => fabric_pd_ready_o(16)
       , fabric_pd_ready_o18                                      => fabric_pd_ready_o(17)
       , fabric_pd_ready_o19                                      => fabric_pd_ready_o(18)
       , fabric_pd_ready_o20                                      => fabric_pd_ready_o(19)
       , fabric_pd_ready_o21                                      => fabric_pd_ready_o(20)
       , fabric_pd_ready_o22                                      => fabric_pd_ready_o(21)
       , fabric_pd_ready_o23                                      => fabric_pd_ready_o(22)
       , fabric_pd_ready_o24                                      => fabric_pd_ready_o(23)
       , fabric_debug_key_correct_o                               => fabric_debug_key_correct_o
       , fabric_otp_apb_ready_o                                   => fabric_otp_apb_ready_o
       , fabric_otp_user_progfail_o                               => fabric_otp_user_progfail_o
       , fabric_mrepair_fuse_sec_o                                => fabric_mrepair_fuse_sec_o
       , fabric_mrepair_fuse_bend2_o                              => fabric_mrepair_fuse_bend2_o
       , fabric_debug_lifecycle_o1                                => fabric_debug_lifecycle_o(0)
       , fabric_debug_lifecycle_o2                                => fabric_debug_lifecycle_o(1)
       , fabric_debug_lifecycle_o3                                => fabric_debug_lifecycle_o(2)
       , fabric_debug_lifecycle_o4                                => fabric_debug_lifecycle_o(3)
       , fabric_mrepair_fuse_ack_o                                => fabric_mrepair_fuse_ack_o
       , fabric_debug_cpt_retry_o1                                => fabric_debug_cpt_retry_o(0)
       , fabric_debug_cpt_retry_o2                                => fabric_debug_cpt_retry_o(1)
       , fabric_debug_cpt_retry_o3                                => fabric_debug_cpt_retry_o(2)
       , fabric_debug_cpt_retry_o4                                => fabric_debug_cpt_retry_o(3)
       , fabric_otp_security_ack_o                                => fabric_otp_security_ack_o
       , fabric_debug_otpmgmt_state_o1                            => fabric_debug_otpmgmt_state_o(0)
       , fabric_debug_otpmgmt_state_o2                            => fabric_debug_otpmgmt_state_o(1)
       , fabric_debug_otpmgmt_state_o3                            => fabric_debug_otpmgmt_state_o(2)
       , fabric_mrepair_fuse_progfail_o                           => fabric_mrepair_fuse_progfail_o
       , fabric_otp_user_bist2fail_o1                             => fabric_otp_user_bist2fail_o(0)
       , fabric_otp_user_bist2fail_o2                             => fabric_otp_user_bist2fail_o(1)
       , fabric_otp_user_bist2fail_o3                             => fabric_otp_user_bist2fail_o(2)
       , fabric_otp_user_bist2fail_o4                             => fabric_otp_user_bist2fail_o(3)
       , fabric_otp_user_bist2fail_o5                             => fabric_otp_user_bist2fail_o(4)
       , fabric_otp_user_bist2fail_o6                             => fabric_otp_user_bist2fail_o(5)
       , fabric_otp_user_bist2fail_o7                             => fabric_otp_user_bist2fail_o(6)
       , fabric_user_data_o1                                      => fabric_user_data_o(0)
       , fabric_user_data_o2                                      => fabric_user_data_o(1)
       , fabric_user_data_o3                                      => fabric_user_data_o(2)
       , fabric_user_data_o4                                      => fabric_user_data_o(3)
       , fabric_user_data_o5                                      => fabric_user_data_o(4)
       , fabric_user_data_o6                                      => fabric_user_data_o(5)
       , fabric_user_data_o7                                      => fabric_user_data_o(6)
       , fabric_user_data_o8                                      => fabric_user_data_o(7)
       , fabric_user_data_o9                                      => fabric_user_data_o(8)
       , fabric_user_data_o10                                     => fabric_user_data_o(9)
       , fabric_user_data_o11                                     => fabric_user_data_o(10)
       , fabric_user_data_o12                                     => fabric_user_data_o(11)
       , fabric_user_data_o13                                     => fabric_user_data_o(12)
       , fabric_user_data_o14                                     => fabric_user_data_o(13)
       , fabric_user_data_o15                                     => fabric_user_data_o(14)
       , fabric_user_data_o16                                     => fabric_user_data_o(15)
       , fabric_user_data_o17                                     => fabric_user_data_o(16)
       , fabric_user_data_o18                                     => fabric_user_data_o(17)
       , fabric_user_data_o19                                     => fabric_user_data_o(18)
       , fabric_user_data_o20                                     => fabric_user_data_o(19)
       , fabric_user_data_o21                                     => fabric_user_data_o(20)
       , fabric_user_data_o22                                     => fabric_user_data_o(21)
       , fabric_user_data_o23                                     => fabric_user_data_o(22)
       , fabric_user_data_o24                                     => fabric_user_data_o(23)
       , fabric_user_data_o25                                     => fabric_user_data_o(24)
       , fabric_user_data_o26                                     => fabric_user_data_o(25)
       , fabric_user_data_o27                                     => fabric_user_data_o(26)
       , fabric_user_data_o28                                     => fabric_user_data_o(27)
       , fabric_user_data_o29                                     => fabric_user_data_o(28)
       , fabric_user_data_o30                                     => fabric_user_data_o(29)
       , fabric_user_data_o31                                     => fabric_user_data_o(30)
       , fabric_user_data_o32                                     => fabric_user_data_o(31)
       , fabric_jtag_tdi_o                                        => fabric_jtag_tdi_o
       , fabric_lowskew_o3                                        => fabric_lowskew_o3
       , fabric_lowskew_o5                                        => fabric_lowskew_o5
       , fabric_lowskew_o4                                        => fabric_lowskew_o4
       , fabric_debug_error_o                                     => fabric_debug_error_o
       , fabric_jtag_usr2_o                                       => fabric_jtag_usr2_o
       , fabric_mrepair_fuse_wlromout_o1                          => fabric_mrepair_fuse_wlromout_o(0)
       , fabric_mrepair_fuse_wlromout_o2                          => fabric_mrepair_fuse_wlromout_o(1)
       , fabric_mrepair_fuse_wlromout_o3                          => fabric_mrepair_fuse_wlromout_o(2)
       , fabric_mrepair_fuse_wlromout_o4                          => fabric_mrepair_fuse_wlromout_o(3)
       , fabric_mrepair_fuse_wlromout_o5                          => fabric_mrepair_fuse_wlromout_o(4)
       , fabric_mrepair_fuse_wlromout_o6                          => fabric_mrepair_fuse_wlromout_o(5)
       , fabric_mrepair_fuse_wlromout_o7                          => fabric_mrepair_fuse_wlromout_o(6)
       , fabric_mrepair_fuse_wlromout_o8                          => fabric_mrepair_fuse_wlromout_o(7)
       , fabric_mrepair_fuse_wlromout_o9                          => fabric_mrepair_fuse_wlromout_o(8)
       , fabric_mrepair_fuse_wlromout_o10                         => fabric_mrepair_fuse_wlromout_o(9)
       , fabric_debug_otpapb_state_o1                             => fabric_debug_otpapb_state_o(0)
       , fabric_debug_otpapb_state_o2                             => fabric_debug_otpapb_state_o(1)
       , fabric_debug_otpapb_state_o3                             => fabric_debug_otpapb_state_o(2)
       , fabric_otp_user_bist1fail_o1                             => fabric_otp_user_bist1fail_o(0)
       , fabric_otp_user_bist1fail_o2                             => fabric_otp_user_bist1fail_o(1)
       , fabric_otp_user_bist1fail_o3                             => fabric_otp_user_bist1fail_o(2)
       , fabric_otp_user_bist1fail_o4                             => fabric_otp_user_bist1fail_o(3)
       , fabric_otp_user_bist1fail_o5                             => fabric_otp_user_bist1fail_o(4)
       , fabric_otp_user_bist1fail_o6                             => fabric_otp_user_bist1fail_o(5)
       , fabric_otp_user_bist1fail_o7                             => fabric_otp_user_bist1fail_o(6)
       , fabric_otp_user_bist1fail_o8                             => fabric_otp_user_bist1fail_o(7)
       , fabric_otp_security_bist_fail2_o1                        => fabric_otp_security_bist_fail2_o(0)
       , fabric_otp_security_bist_fail2_o2                        => fabric_otp_security_bist_fail2_o(1)
       , fabric_otp_security_bist_fail2_o3                        => fabric_otp_security_bist_fail2_o(2)
       , fabric_otp_security_bist_fail2_o4                        => fabric_otp_security_bist_fail2_o(3)
       , fabric_otp_security_bist_fail2_o5                        => fabric_otp_security_bist_fail2_o(4)
       , fabric_otp_security_bist_fail2_o6                        => fabric_otp_security_bist_fail2_o(5)
       , fabric_otp_security_bist_fail2_o7                        => fabric_otp_security_bist_fail2_o(6)
       , fabric_otp_user_disturbed_o                              => fabric_otp_user_disturbed_o
       , fabric_flag_trigger_o                                    => fabric_flag_trigger_o
       , fabric_otp_security_bist_end2_o                          => fabric_otp_security_bist_end2_o
       , fabric_otp_security_bist_fail1_o1                        => fabric_otp_security_bist_fail1_o(0)
       , fabric_otp_security_bist_fail1_o2                        => fabric_otp_security_bist_fail1_o(1)
       , fabric_otp_security_bist_fail1_o3                        => fabric_otp_security_bist_fail1_o(2)
       , fabric_otp_security_bist_fail1_o4                        => fabric_otp_security_bist_fail1_o(3)
       , fabric_otp_security_bist_fail1_o5                        => fabric_otp_security_bist_fail1_o(4)
       , fabric_otp_security_bist_fail1_o6                        => fabric_otp_security_bist_fail1_o(5)
       , fabric_otp_security_bist_fail1_o7                        => fabric_otp_security_bist_fail1_o(6)
       , fabric_otp_security_bist_fail1_o8                        => fabric_otp_security_bist_fail1_o(7)
       , fabric_mrepair_fuse_locked_o                             => fabric_mrepair_fuse_locked_o
       , fabric_otp_user_flagstate_o1                             => fabric_otp_user_flagstate_o(0)
       , fabric_otp_user_flagstate_o2                             => fabric_otp_user_flagstate_o(1)
       , fabric_otp_user_flagstate_o3                             => fabric_otp_user_flagstate_o(2)
       , fabric_otp_user_flagstate_o4                             => fabric_otp_user_flagstate_o(3)
       , fabric_otp_security_scanout_o1                           => fabric_otp_security_scanout_o(0)
       , fabric_otp_security_scanout_o2                           => fabric_otp_security_scanout_o(1)
       , fabric_otp_security_scanout_o3                           => fabric_otp_security_scanout_o(2)
       , fabric_otp_security_scanout_o4                           => fabric_otp_security_scanout_o(3)
       , fabric_otp_security_scanout_o5                           => fabric_otp_security_scanout_o(4)
       , fabric_user_write_cycle_o                                => fabric_user_write_cycle_o
       , fabric_debug_fsm_state_o1                                => fabric_debug_fsm_state_o(0)
       , fabric_debug_fsm_state_o2                                => fabric_debug_fsm_state_o(1)
       , fabric_debug_fsm_state_o3                                => fabric_debug_fsm_state_o(2)
       , fabric_otp_user_ded_o                                    => fabric_otp_user_ded_o
       , fabric_debug_otp_manager_read_done_o                     => fabric_debug_otp_manager_read_done_o
       , fabric_debug_frame_use_encryption_o                      => fabric_debug_frame_use_encryption_o
       , fabric_data_to_system_o                                  => fabric_data_to_system_o
       , fabric_jtag_usr1_o                                       => fabric_jtag_usr1_o
       , fabric_otp_user_bend1_o                                  => fabric_otp_user_bend1_o
       , fabric_debug_otpboot_curr_addr_o1                        => fabric_debug_otpboot_curr_addr_o(0)
       , fabric_debug_otpboot_curr_addr_o2                        => fabric_debug_otpboot_curr_addr_o(1)
       , fabric_debug_otpboot_curr_addr_o3                        => fabric_debug_otpboot_curr_addr_o(2)
       , fabric_debug_otpboot_curr_addr_o4                        => fabric_debug_otpboot_curr_addr_o(3)
       , fabric_debug_otpboot_curr_addr_o5                        => fabric_debug_otpboot_curr_addr_o(4)
       , fabric_debug_otpboot_curr_addr_o6                        => fabric_debug_otpboot_curr_addr_o(5)
       , fabric_debug_otpboot_curr_addr_o7                        => fabric_debug_otpboot_curr_addr_o(6)
       , fabric_debug_otpboot_curr_addr_o8                        => fabric_debug_otpboot_curr_addr_o(7)
       , fabric_mrepair_fuse_ready_o                              => fabric_mrepair_fuse_ready_o
       , fabric_mrepair_fuse_calibrated_o                         => fabric_mrepair_fuse_calibrated_o
       , fabric_sif_load_en_to_bist_o1                            => fabric_sif_load_en_to_bist_o(0)
       , fabric_sif_load_en_to_bist_o2                            => fabric_sif_load_en_to_bist_o(1)
       , fabric_sif_load_en_to_bist_o3                            => fabric_sif_load_en_to_bist_o(2)
       , fabric_sif_load_en_to_bist_o4                            => fabric_sif_load_en_to_bist_o(3)
       , fabric_sif_load_en_to_bist_o5                            => fabric_sif_load_en_to_bist_o(4)
       , fabric_sif_load_en_to_bist_o6                            => fabric_sif_load_en_to_bist_o(5)
       , fabric_sif_load_en_to_bist_o7                            => fabric_sif_load_en_to_bist_o(6)
       , fabric_sif_load_en_to_bist_o8                            => fabric_sif_load_en_to_bist_o(7)
       , fabric_sif_load_en_to_bist_o9                            => fabric_sif_load_en_to_bist_o(8)
       , fabric_sif_load_en_to_bist_o10                           => fabric_sif_load_en_to_bist_o(9)
       , fabric_sif_load_en_to_bist_o11                           => fabric_sif_load_en_to_bist_o(10)
       , fabric_sif_load_en_to_bist_o12                           => fabric_sif_load_en_to_bist_o(11)
       , fabric_sif_load_en_to_bist_o13                           => fabric_sif_load_en_to_bist_o(12)
       , fabric_sif_load_en_to_bist_o14                           => fabric_sif_load_en_to_bist_o(13)
       , fabric_sif_load_en_to_bist_o15                           => fabric_sif_load_en_to_bist_o(14)
       , fabric_sif_load_en_to_bist_o16                           => fabric_sif_load_en_to_bist_o(15)
       , fabric_sif_load_en_to_bist_o17                           => fabric_sif_load_en_to_bist_o(16)
       , fabric_sif_load_en_to_bist_o18                           => fabric_sif_load_en_to_bist_o(17)
       , fabric_sif_load_en_to_bist_o19                           => fabric_sif_load_en_to_bist_o(18)
       , fabric_sif_load_en_to_bist_o20                           => fabric_sif_load_en_to_bist_o(19)
       , fabric_sif_load_en_to_bist_o21                           => fabric_sif_load_en_to_bist_o(20)
       , fabric_sif_load_en_to_bist_o22                           => fabric_sif_load_en_to_bist_o(21)
       , fabric_sif_load_en_to_bist_o23                           => fabric_sif_load_en_to_bist_o(22)
       , fabric_sif_load_en_to_bist_o24                           => fabric_sif_load_en_to_bist_o(23)
       , fabric_io_out_o1                                         => fabric_io_out_o(0)
       , fabric_io_out_o2                                         => fabric_io_out_o(1)
       , fabric_io_out_o3                                         => fabric_io_out_o(2)
       , fabric_io_out_o4                                         => fabric_io_out_o(3)
       , fabric_io_out_o5                                         => fabric_io_out_o(4)
       , fabric_io_out_o6                                         => fabric_io_out_o(5)
       , fabric_io_out_o7                                         => fabric_io_out_o(6)
       , fabric_io_out_o8                                         => fabric_io_out_o(7)
       , fabric_io_out_o9                                         => fabric_io_out_o(8)
       , fabric_io_out_o10                                        => fabric_io_out_o(9)
       , fabric_io_out_o11                                        => fabric_io_out_o(10)
       , fabric_io_out_o12                                        => fabric_io_out_o(11)
       , fabric_io_out_o13                                        => fabric_io_out_o(12)
       , fabric_io_out_o14                                        => fabric_io_out_o(13)
       , fabric_io_out_o15                                        => fabric_io_out_o(14)
       , fabric_io_out_o16                                        => fabric_io_out_o(15)
       , fabric_io_out_o17                                        => fabric_io_out_o(16)
       , fabric_io_out_o18                                        => fabric_io_out_o(17)
       , fabric_io_out_o19                                        => fabric_io_out_o(18)
       , fabric_io_out_o20                                        => fabric_io_out_o(19)
       , fabric_io_out_o21                                        => fabric_io_out_o(20)
       , fabric_io_out_o22                                        => fabric_io_out_o(21)
       , fabric_io_out_o23                                        => fabric_io_out_o(22)
       , fabric_io_out_o24                                        => fabric_io_out_o(23)
       , fabric_io_out_o25                                        => fabric_io_out_o(24)
       , fabric_mrepair_fuse_startword_o1                         => fabric_mrepair_fuse_startword_o(0)
       , fabric_mrepair_fuse_startword_o2                         => fabric_mrepair_fuse_startword_o(1)
       , fabric_mrepair_fuse_startword_o3                         => fabric_mrepair_fuse_startword_o(2)
       , fabric_mrepair_fuse_startword_o4                         => fabric_mrepair_fuse_startword_o(3)
       , fabric_mrepair_fuse_startword_o5                         => fabric_mrepair_fuse_startword_o(4)
       , fabric_mrepair_fuse_startword_o6                         => fabric_mrepair_fuse_startword_o(5)
       , fabric_mrepair_fuse_startword_o7                         => fabric_mrepair_fuse_startword_o(6)
       , fabric_mrepair_fuse_startword_o8                         => fabric_mrepair_fuse_startword_o(7)
       , fabric_mrepair_fuse_startword_o9                         => fabric_mrepair_fuse_startword_o(8)
       , fabric_mrepair_fuse_startword_o10                        => fabric_mrepair_fuse_startword_o(9)
       , fabric_mrepair_fuse_startword_o11                        => fabric_mrepair_fuse_startword_o(10)
       , fabric_mrepair_fuse_startword_o12                        => fabric_mrepair_fuse_startword_o(11)
       , fabric_mrepair_fuse_startword_o13                        => fabric_mrepair_fuse_startword_o(12)
       , fabric_mrepair_fuse_startword_o14                        => fabric_mrepair_fuse_startword_o(13)
       , fabric_mrepair_fuse_startword_o15                        => fabric_mrepair_fuse_startword_o(14)
       , fabric_mrepair_fuse_startword_o16                        => fabric_mrepair_fuse_startword_o(15)
       , fabric_system_dataready_o                                => fabric_system_dataready_o
       , fabric_mrepair_fuse_pwok_o                               => fabric_mrepair_fuse_pwok_o
       , fabric_lowskew_o6                                        => fabric_lowskew_o6
       , fabric_cfg_fabric_user_flag_o                            => fabric_cfg_fabric_user_flag_o
       , fabric_otp_user_dout_o1                                  => fabric_otp_user_dout_o(0)
       , fabric_otp_user_dout_o2                                  => fabric_otp_user_dout_o(1)
       , fabric_otp_user_dout_o3                                  => fabric_otp_user_dout_o(2)
       , fabric_otp_user_dout_o4                                  => fabric_otp_user_dout_o(3)
       , fabric_otp_user_dout_o5                                  => fabric_otp_user_dout_o(4)
       , fabric_otp_user_dout_o6                                  => fabric_otp_user_dout_o(5)
       , fabric_otp_user_dout_o7                                  => fabric_otp_user_dout_o(6)
       , fabric_otp_user_dout_o8                                  => fabric_otp_user_dout_o(7)
       , fabric_otp_user_dout_o9                                  => fabric_otp_user_dout_o(8)
       , fabric_otp_user_dout_o10                                 => fabric_otp_user_dout_o(9)
       , fabric_otp_user_dout_o11                                 => fabric_otp_user_dout_o(10)
       , fabric_otp_user_dout_o12                                 => fabric_otp_user_dout_o(11)
       , fabric_otp_user_dout_o13                                 => fabric_otp_user_dout_o(12)
       , fabric_otp_user_dout_o14                                 => fabric_otp_user_dout_o(13)
       , fabric_otp_user_dout_o15                                 => fabric_otp_user_dout_o(14)
       , fabric_otp_user_dout_o16                                 => fabric_otp_user_dout_o(15)
       , fabric_otp_user_dout_o17                                 => fabric_otp_user_dout_o(16)
       , fabric_otp_user_dout_o18                                 => fabric_otp_user_dout_o(17)
       , fabric_otp_user_dout_o19                                 => fabric_otp_user_dout_o(18)
       , fabric_otp_user_dout_o20                                 => fabric_otp_user_dout_o(19)
       , fabric_otp_user_dout_o21                                 => fabric_otp_user_dout_o(20)
       , fabric_otp_user_dout_o22                                 => fabric_otp_user_dout_o(21)
       , fabric_otp_user_dout_o23                                 => fabric_otp_user_dout_o(22)
       , fabric_otp_user_dout_o24                                 => fabric_otp_user_dout_o(23)
       , fabric_otp_user_dout_o25                                 => fabric_otp_user_dout_o(24)
       , fabric_otp_user_dout_o26                                 => fabric_otp_user_dout_o(25)
       , fabric_otp_user_dout_o27                                 => fabric_otp_user_dout_o(26)
       , fabric_otp_user_dout_o28                                 => fabric_otp_user_dout_o(27)
       , fabric_otp_user_dout_o29                                 => fabric_otp_user_dout_o(28)
       , fabric_otp_user_dout_o30                                 => fabric_otp_user_dout_o(29)
       , fabric_otp_user_dout_o31                                 => fabric_otp_user_dout_o(30)
       , fabric_otp_user_dout_o32                                 => fabric_otp_user_dout_o(31)
       , fabric_otp_user_dout_o33                                 => fabric_otp_user_dout_o(32)
       , fabric_otp_user_dout_o34                                 => fabric_otp_user_dout_o(33)
       , fabric_otp_user_dout_o35                                 => fabric_otp_user_dout_o(34)
       , fabric_otp_user_dout_o36                                 => fabric_otp_user_dout_o(35)
       , fabric_otp_user_dout_o37                                 => fabric_otp_user_dout_o(36)
       , fabric_otp_user_dout_o38                                 => fabric_otp_user_dout_o(37)
       , fabric_otp_user_dout_o39                                 => fabric_otp_user_dout_o(38)
       , fabric_otp_user_dout_o40                                 => fabric_otp_user_dout_o(39)
       , fabric_otp_user_dout_o41                                 => fabric_otp_user_dout_o(40)
       , fabric_mrepair_fuse_bist2fail_o1                         => fabric_mrepair_fuse_bist2fail_o(0)
       , fabric_mrepair_fuse_bist2fail_o2                         => fabric_mrepair_fuse_bist2fail_o(1)
       , fabric_mrepair_fuse_bist2fail_o3                         => fabric_mrepair_fuse_bist2fail_o(2)
       , fabric_mrepair_fuse_bist2fail_o4                         => fabric_mrepair_fuse_bist2fail_o(3)
       , fabric_mrepair_fuse_bist2fail_o5                         => fabric_mrepair_fuse_bist2fail_o(4)
       , fabric_mrepair_fuse_bist2fail_o6                         => fabric_mrepair_fuse_bist2fail_o(5)
       , fabric_mrepair_fuse_bist2fail_o7                         => fabric_mrepair_fuse_bist2fail_o(6)
       , fabric_status_cold_start_o                               => fabric_status_cold_start_o
       , fabric_flag_error_o                                      => fabric_flag_error_o
       , fabric_debug_direct_permission_read_o1                   => fabric_debug_direct_permission_read_o(0)
       , fabric_debug_direct_permission_read_o2                   => fabric_debug_direct_permission_read_o(1)
       , fabric_debug_direct_permission_read_o3                   => fabric_debug_direct_permission_read_o(2)
       , fabric_debug_direct_permission_read_o4                   => fabric_debug_direct_permission_read_o(3)
);
end NX_ARCH;
-- =================================================================================================
--  NX_SOC_INTERFACE definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_SOC_INTERFACE is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    -- dahlia <-> fabric
    fabric_lowskew_o1                            : out std_logic;  -- dahlia_clk_fpga_i
    fabric_lowskew_i1                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i2                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i3                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i4                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i5                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i6                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i7                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i8                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i9                            : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_i10                           : in  std_logic;  -- dahlia_clk_fpga_nic_o
    fabric_lowskew_o2                            : out std_logic;  -- dahlia_rstn_fpga_out_i
    fabric_fpga_nic_rstn_i1                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i2                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i3                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i4                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i5                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i6                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i7                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i8                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i9                      : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_nic_rstn_i10                     : in  std_logic;  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_pmrstn_i                         : in  std_logic;  -- dahlia_fpga_pmrstn_o
    fabric_fpga_sysrstn_i                        : in  std_logic;  -- dahlia_fpga_sysrstn_o
    fabric_fpga_trigger_in_o1                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o2                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o3                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o4                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o5                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o6                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o7                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_in_o8                    : out std_logic;  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_out_i1                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i2                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i3                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i4                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i5                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i6                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i7                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_trigger_out_i8                   : in  std_logic;  -- dahlia_fpga_trigger_out_o
    fabric_fpga_interrupt_in_i1                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i2                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i3                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i4                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i5                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i6                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i7                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i8                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i9                  : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i10                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i11                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i12                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i13                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i14                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i15                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i16                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i17                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i18                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i19                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i20                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i21                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i22                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i23                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i24                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i25                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i26                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i27                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i28                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i29                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i30                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i31                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i32                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i33                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i34                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i35                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i36                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i37                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i38                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i39                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i40                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i41                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i42                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i43                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i44                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i45                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i46                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i47                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i48                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i49                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i50                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i51                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i52                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i53                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i54                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i55                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i56                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i57                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i58                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i59                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i60                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i61                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i62                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i63                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i64                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i65                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i66                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i67                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i68                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i69                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i70                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i71                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i72                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i73                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i74                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i75                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i76                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i77                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i78                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i79                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i80                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i81                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i82                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i83                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i84                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i85                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i86                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i87                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i88                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i89                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i90                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i91                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i92                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i93                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i94                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i95                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i96                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i97                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i98                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i99                 : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i100                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i101                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i102                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i103                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i104                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i105                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i106                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i107                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i108                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i109                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i110                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i111                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i112                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i113                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i114                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i115                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i116                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i117                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i118                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i119                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_fpga_interrupt_in_i120                : in  std_logic;  -- dahlia_fpga_interrupt_in_o
    fabric_sysc_hold_on_debug_i                  : in  std_logic;  -- dahlia_sysc_hold_on_debug_o
    fabric_fpga_events60_i1                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i2                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i3                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i4                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i5                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i6                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i7                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i8                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i9                      : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i10                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i11                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i12                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i13                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i14                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i15                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i16                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i17                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i18                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i19                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i20                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i21                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i22                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i23                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i24                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i25                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i26                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i27                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i28                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i29                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i30                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i31                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i32                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i33                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i34                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i35                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i36                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i37                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i38                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i39                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i40                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i41                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i42                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i43                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i44                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i45                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i46                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i47                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i48                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i49                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i50                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i51                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i52                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i53                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i54                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i55                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i56                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i57                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i58                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i59                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_events60_i60                     : in  std_logic;  -- dahlia_fpga_events60_o
    fabric_fpga_araddr_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o4                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o5                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o6                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o7                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o8                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o9                 : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o10                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o11                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o12                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o13                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o14                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o15                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o16                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o17                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o18                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o19                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o20                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o21                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o22                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o23                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o24                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o25                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o26                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o27                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o28                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o29                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o30                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o31                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o32                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o33                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o34                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o35                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o36                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o37                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o38                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o39                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_araddr_axi_s1_o40                : out std_logic;  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_arburst_axi_s1_o1                : out std_logic;  -- dahlia_fpga_arburst_axi_s1_i
    fabric_fpga_arburst_axi_s1_o2                : out std_logic;  -- dahlia_fpga_arburst_axi_s1_i
    fabric_fpga_arcache_axi_s1_o1                : out std_logic;  -- dahlia_fpga_arcache_axi_s1_i
    fabric_fpga_arcache_axi_s1_o2                : out std_logic;  -- dahlia_fpga_arcache_axi_s1_i
    fabric_fpga_arcache_axi_s1_o3                : out std_logic;  -- dahlia_fpga_arcache_axi_s1_i
    fabric_fpga_arcache_axi_s1_o4                : out std_logic;  -- dahlia_fpga_arcache_axi_s1_i
    fabric_fpga_arid_axi_s1_o1                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o2                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o3                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o4                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o5                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o6                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o7                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o8                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o9                   : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o10                  : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o11                  : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arid_axi_s1_o12                  : out std_logic;  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arlen_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o5                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o6                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o7                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlen_axi_s1_o8                  : out std_logic;  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlock_axi_s1_o                  : out std_logic;  -- dahlia_fpga_arlock_axi_s1_i
    fabric_fpga_arprot_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_arprot_axi_s1_i
    fabric_fpga_arprot_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_arprot_axi_s1_i
    fabric_fpga_arprot_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_arprot_axi_s1_i
    fabric_fpga_arqos_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_arqos_axi_s1_i
    fabric_fpga_arqos_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_arqos_axi_s1_i
    fabric_fpga_arqos_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_arqos_axi_s1_i
    fabric_fpga_arqos_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_arqos_axi_s1_i
    fabric_fpga_arregion_axi_s1_o1               : out std_logic;  -- dahlia_fpga_arregion_axi_s1_i
    fabric_fpga_arregion_axi_s1_o2               : out std_logic;  -- dahlia_fpga_arregion_axi_s1_i
    fabric_fpga_arregion_axi_s1_o3               : out std_logic;  -- dahlia_fpga_arregion_axi_s1_i
    fabric_fpga_arregion_axi_s1_o4               : out std_logic;  -- dahlia_fpga_arregion_axi_s1_i
    fabric_fpga_arsize_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_arsize_axi_s1_i
    fabric_fpga_arsize_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_arsize_axi_s1_i
    fabric_fpga_arsize_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_arsize_axi_s1_i
    fabric_fpga_arvalid_axi_s1_o                 : out std_logic;  -- dahlia_fpga_arvalid_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o4                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o5                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o6                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o7                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o8                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o9                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o10                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o11                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o12                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o13                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o14                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o15                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o16                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o17                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o18                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o19                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o20                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o21                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o22                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o23                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o24                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o25                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o26                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o27                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o28                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o29                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o30                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o31                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o32                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o33                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o34                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o35                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o36                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o37                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o38                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o39                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o40                : out std_logic;  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awburst_axi_s1_o1                : out std_logic;  -- dahlia_fpga_awburst_axi_s1_i
    fabric_fpga_awburst_axi_s1_o2                : out std_logic;  -- dahlia_fpga_awburst_axi_s1_i
    fabric_fpga_awcache_axi_s1_o1                : out std_logic;  -- dahlia_fpga_awcache_axi_s1_i
    fabric_fpga_awcache_axi_s1_o2                : out std_logic;  -- dahlia_fpga_awcache_axi_s1_i
    fabric_fpga_awcache_axi_s1_o3                : out std_logic;  -- dahlia_fpga_awcache_axi_s1_i
    fabric_fpga_awcache_axi_s1_o4                : out std_logic;  -- dahlia_fpga_awcache_axi_s1_i
    fabric_fpga_awid_axi_s1_o1                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o2                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o3                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o4                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o5                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o6                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o7                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o8                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o9                   : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o10                  : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o11                  : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awid_axi_s1_o12                  : out std_logic;  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awlen_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o5                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o6                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o7                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlen_axi_s1_o8                  : out std_logic;  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlock_axi_s1_o                  : out std_logic;  -- dahlia_fpga_awlock_axi_s1_i
    fabric_fpga_awprot_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_awprot_axi_s1_i
    fabric_fpga_awprot_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_awprot_axi_s1_i
    fabric_fpga_awprot_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_awprot_axi_s1_i
    fabric_fpga_awqos_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_awqos_axi_s1_i
    fabric_fpga_awqos_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_awqos_axi_s1_i
    fabric_fpga_awqos_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_awqos_axi_s1_i
    fabric_fpga_awqos_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_awqos_axi_s1_i
    fabric_fpga_awregion_axi_s1_o1               : out std_logic;  -- dahlia_fpga_awregion_axi_s1_i
    fabric_fpga_awregion_axi_s1_o2               : out std_logic;  -- dahlia_fpga_awregion_axi_s1_i
    fabric_fpga_awregion_axi_s1_o3               : out std_logic;  -- dahlia_fpga_awregion_axi_s1_i
    fabric_fpga_awregion_axi_s1_o4               : out std_logic;  -- dahlia_fpga_awregion_axi_s1_i
    fabric_fpga_awsize_axi_s1_o1                 : out std_logic;  -- dahlia_fpga_awsize_axi_s1_i
    fabric_fpga_awsize_axi_s1_o2                 : out std_logic;  -- dahlia_fpga_awsize_axi_s1_i
    fabric_fpga_awsize_axi_s1_o3                 : out std_logic;  -- dahlia_fpga_awsize_axi_s1_i
    fabric_fpga_bready_axi_s1_o                  : out std_logic;  -- dahlia_fpga_bready_axi_s1_i
    fabric_fpga_rready_axi_s1_o                  : out std_logic;  -- dahlia_fpga_rready_axi_s1_i
    fabric_fpga_wdata_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o5                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o6                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o7                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o8                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o9                  : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o10                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o11                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o12                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o13                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o14                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o15                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o16                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o17                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o18                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o19                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o20                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o21                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o22                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o23                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o24                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o25                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o26                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o27                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o28                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o29                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o30                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o31                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o32                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o33                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o34                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o35                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o36                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o37                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o38                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o39                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o40                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o41                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o42                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o43                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o44                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o45                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o46                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o47                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o48                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o49                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o50                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o51                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o52                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o53                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o54                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o55                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o56                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o57                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o58                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o59                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o60                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o61                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o62                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o63                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o64                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o65                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o66                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o67                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o68                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o69                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o70                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o71                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o72                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o73                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o74                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o75                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o76                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o77                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o78                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o79                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o80                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o81                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o82                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o83                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o84                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o85                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o86                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o87                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o88                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o89                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o90                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o91                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o92                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o93                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o94                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o95                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o96                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o97                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o98                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o99                 : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o100                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o101                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o102                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o103                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o104                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o105                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o106                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o107                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o108                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o109                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o110                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o111                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o112                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o113                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o114                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o115                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o116                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o117                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o118                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o119                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o120                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o121                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o122                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o123                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o124                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o125                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o126                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o127                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wdata_axi_s1_o128                : out std_logic;  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wlast_axi_s1_o                   : out std_logic;  -- dahlia_fpga_wlast_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o1                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o2                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o3                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o4                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o5                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o6                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o7                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o8                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o9                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o10                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o11                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o12                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o13                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o14                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o15                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o16                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wvalid_axi_s1_o                  : out std_logic;  -- dahlia_fpga_wvalid_axi_s1_i
    fabric_fpga_awvalid_axi_s1_o                 : out std_logic;  -- dahlia_fpga_awvalid_axi_s1_i
    fabric_fpga_arready_axi_s1_i                 : in  std_logic;  -- dahlia_fpga_arready_axi_s1_o
    fabric_fpga_awready_axi_s1_i                 : in  std_logic;  -- dahlia_fpga_awready_axi_s1_o
    fabric_fpga_bid_axi_s1_i1                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i2                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i3                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i4                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i5                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i6                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i7                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i8                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i9                    : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i10                   : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i11                   : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bid_axi_s1_i12                   : in  std_logic;  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bresp_axi_s1_i1                  : in  std_logic;  -- dahlia_fpga_bresp_axi_s1_o
    fabric_fpga_bresp_axi_s1_i2                  : in  std_logic;  -- dahlia_fpga_bresp_axi_s1_o
    fabric_fpga_bvalid_axi_s1_i                  : in  std_logic;  -- dahlia_fpga_bvalid_axi_s1_o
    fabric_fpga_rdata_axi_s1_i1                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i2                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i3                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i4                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i5                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i6                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i7                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i8                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i9                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i10                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i11                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i12                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i13                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i14                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i15                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i16                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i17                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i18                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i19                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i20                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i21                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i22                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i23                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i24                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i25                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i26                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i27                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i28                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i29                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i30                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i31                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i32                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i33                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i34                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i35                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i36                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i37                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i38                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i39                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i40                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i41                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i42                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i43                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i44                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i45                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i46                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i47                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i48                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i49                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i50                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i51                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i52                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i53                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i54                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i55                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i56                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i57                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i58                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i59                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i60                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i61                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i62                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i63                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i64                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i65                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i66                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i67                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i68                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i69                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i70                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i71                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i72                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i73                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i74                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i75                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i76                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i77                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i78                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i79                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i80                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i81                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i82                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i83                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i84                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i85                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i86                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i87                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i88                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i89                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i90                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i91                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i92                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i93                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i94                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i95                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i96                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i97                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i98                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i99                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i100                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i101                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i102                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i103                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i104                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i105                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i106                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i107                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i108                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i109                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i110                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i111                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i112                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i113                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i114                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i115                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i116                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i117                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i118                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i119                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i120                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i121                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i122                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i123                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i124                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i125                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i126                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i127                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rdata_axi_s1_i128                : in  std_logic;  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rid_axi_s1_i1                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i2                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i3                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i4                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i5                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i6                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i7                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i8                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i9                    : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i10                   : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i11                   : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rid_axi_s1_i12                   : in  std_logic;  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rlast_axi_s1_i                   : in  std_logic;  -- dahlia_fpga_rlast_axi_s1_o
    fabric_fpga_rresp_axi_s1_i1                  : in  std_logic;  -- dahlia_fpga_rresp_axi_s1_o
    fabric_fpga_rresp_axi_s1_i2                  : in  std_logic;  -- dahlia_fpga_rresp_axi_s1_o
    fabric_fpga_rvalid_axi_s1_i                  : in  std_logic;  -- dahlia_fpga_rvalid_axi_s1_o
    fabric_fpga_wready_axi_s1_i                  : in  std_logic;  -- dahlia_fpga_wready_axi_s1_o
    fabric_fpga_araddr_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o4                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o5                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o6                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o7                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o8                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o9                 : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o10                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o11                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o12                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o13                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o14                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o15                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o16                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o17                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o18                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o19                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o20                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o21                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o22                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o23                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o24                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o25                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o26                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o27                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o28                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o29                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o30                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o31                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o32                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o33                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o34                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o35                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o36                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o37                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o38                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o39                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_araddr_axi_s2_o40                : out std_logic;  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_arburst_axi_s2_o1                : out std_logic;  -- dahlia_fpga_arburst_axi_s2_i
    fabric_fpga_arburst_axi_s2_o2                : out std_logic;  -- dahlia_fpga_arburst_axi_s2_i
    fabric_fpga_arcache_axi_s2_o1                : out std_logic;  -- dahlia_fpga_arcache_axi_s2_i
    fabric_fpga_arcache_axi_s2_o2                : out std_logic;  -- dahlia_fpga_arcache_axi_s2_i
    fabric_fpga_arcache_axi_s2_o3                : out std_logic;  -- dahlia_fpga_arcache_axi_s2_i
    fabric_fpga_arcache_axi_s2_o4                : out std_logic;  -- dahlia_fpga_arcache_axi_s2_i
    fabric_fpga_arid_axi_s2_o1                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o2                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o3                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o4                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o5                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o6                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o7                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o8                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o9                   : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o10                  : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o11                  : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arid_axi_s2_o12                  : out std_logic;  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arlen_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o5                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o6                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o7                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlen_axi_s2_o8                  : out std_logic;  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlock_axi_s2_o                  : out std_logic;  -- dahlia_fpga_arlock_axi_s2_i
    fabric_fpga_arprot_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_arprot_axi_s2_i
    fabric_fpga_arprot_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_arprot_axi_s2_i
    fabric_fpga_arprot_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_arprot_axi_s2_i
    fabric_fpga_arqos_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_arqos_axi_s2_i
    fabric_fpga_arqos_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_arqos_axi_s2_i
    fabric_fpga_arqos_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_arqos_axi_s2_i
    fabric_fpga_arqos_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_arqos_axi_s2_i
    fabric_fpga_arregion_axi_s2_o1               : out std_logic;  -- dahlia_fpga_arregion_axi_s2_i
    fabric_fpga_arregion_axi_s2_o2               : out std_logic;  -- dahlia_fpga_arregion_axi_s2_i
    fabric_fpga_arregion_axi_s2_o3               : out std_logic;  -- dahlia_fpga_arregion_axi_s2_i
    fabric_fpga_arregion_axi_s2_o4               : out std_logic;  -- dahlia_fpga_arregion_axi_s2_i
    fabric_fpga_arsize_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_arsize_axi_s2_i
    fabric_fpga_arsize_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_arsize_axi_s2_i
    fabric_fpga_arsize_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_arsize_axi_s2_i
    fabric_fpga_arvalid_axi_s2_o                 : out std_logic;  -- dahlia_fpga_arvalid_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o4                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o5                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o6                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o7                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o8                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o9                 : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o10                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o11                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o12                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o13                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o14                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o15                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o16                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o17                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o18                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o19                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o20                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o21                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o22                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o23                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o24                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o25                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o26                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o27                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o28                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o29                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o30                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o31                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o32                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o33                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o34                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o35                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o36                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o37                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o38                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o39                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o40                : out std_logic;  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awburst_axi_s2_o1                : out std_logic;  -- dahlia_fpga_awburst_axi_s2_i
    fabric_fpga_awburst_axi_s2_o2                : out std_logic;  -- dahlia_fpga_awburst_axi_s2_i
    fabric_fpga_awcache_axi_s2_o1                : out std_logic;  -- dahlia_fpga_awcache_axi_s2_i
    fabric_fpga_awcache_axi_s2_o2                : out std_logic;  -- dahlia_fpga_awcache_axi_s2_i
    fabric_fpga_awcache_axi_s2_o3                : out std_logic;  -- dahlia_fpga_awcache_axi_s2_i
    fabric_fpga_awcache_axi_s2_o4                : out std_logic;  -- dahlia_fpga_awcache_axi_s2_i
    fabric_fpga_awid_axi_s2_o1                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o2                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o3                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o4                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o5                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o6                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o7                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o8                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o9                   : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o10                  : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o11                  : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awid_axi_s2_o12                  : out std_logic;  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awlen_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o5                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o6                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o7                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlen_axi_s2_o8                  : out std_logic;  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlock_axi_s2_o                  : out std_logic;  -- dahlia_fpga_awlock_axi_s2_i
    fabric_fpga_awprot_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_awprot_axi_s2_i
    fabric_fpga_awprot_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_awprot_axi_s2_i
    fabric_fpga_awprot_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_awprot_axi_s2_i
    fabric_fpga_awqos_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_awqos_axi_s2_i
    fabric_fpga_awqos_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_awqos_axi_s2_i
    fabric_fpga_awqos_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_awqos_axi_s2_i
    fabric_fpga_awqos_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_awqos_axi_s2_i
    fabric_fpga_awregion_axi_s2_o1               : out std_logic;  -- dahlia_fpga_awregion_axi_s2_i
    fabric_fpga_awregion_axi_s2_o2               : out std_logic;  -- dahlia_fpga_awregion_axi_s2_i
    fabric_fpga_awregion_axi_s2_o3               : out std_logic;  -- dahlia_fpga_awregion_axi_s2_i
    fabric_fpga_awregion_axi_s2_o4               : out std_logic;  -- dahlia_fpga_awregion_axi_s2_i
    fabric_fpga_awsize_axi_s2_o1                 : out std_logic;  -- dahlia_fpga_awsize_axi_s2_i
    fabric_fpga_awsize_axi_s2_o2                 : out std_logic;  -- dahlia_fpga_awsize_axi_s2_i
    fabric_fpga_awsize_axi_s2_o3                 : out std_logic;  -- dahlia_fpga_awsize_axi_s2_i
    fabric_fpga_bready_axi_s2_o                  : out std_logic;  -- dahlia_fpga_bready_axi_s2_i
    fabric_fpga_rready_axi_s2_o                  : out std_logic;  -- dahlia_fpga_rready_axi_s2_i
    fabric_fpga_wdata_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o5                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o6                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o7                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o8                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o9                  : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o10                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o11                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o12                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o13                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o14                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o15                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o16                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o17                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o18                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o19                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o20                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o21                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o22                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o23                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o24                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o25                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o26                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o27                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o28                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o29                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o30                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o31                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o32                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o33                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o34                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o35                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o36                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o37                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o38                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o39                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o40                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o41                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o42                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o43                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o44                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o45                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o46                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o47                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o48                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o49                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o50                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o51                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o52                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o53                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o54                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o55                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o56                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o57                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o58                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o59                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o60                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o61                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o62                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o63                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o64                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o65                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o66                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o67                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o68                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o69                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o70                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o71                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o72                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o73                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o74                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o75                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o76                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o77                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o78                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o79                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o80                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o81                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o82                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o83                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o84                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o85                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o86                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o87                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o88                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o89                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o90                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o91                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o92                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o93                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o94                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o95                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o96                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o97                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o98                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o99                 : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o100                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o101                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o102                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o103                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o104                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o105                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o106                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o107                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o108                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o109                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o110                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o111                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o112                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o113                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o114                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o115                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o116                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o117                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o118                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o119                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o120                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o121                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o122                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o123                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o124                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o125                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o126                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o127                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wdata_axi_s2_o128                : out std_logic;  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wlast_axi_s2_o                   : out std_logic;  -- dahlia_fpga_wlast_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o1                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o2                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o3                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o4                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o5                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o6                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o7                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o8                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o9                  : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o10                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o11                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o12                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o13                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o14                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o15                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o16                 : out std_logic;  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wvalid_axi_s2_o                  : out std_logic;  -- dahlia_fpga_wvalid_axi_s2_i
    fabric_fpga_awvalid_axi_s2_o                 : out std_logic;  -- dahlia_fpga_awvalid_axi_s2_i
    fabric_fpga_arready_axi_s2_i                 : in  std_logic;  -- dahlia_fpga_arready_axi_s2_o
    fabric_fpga_awready_axi_s2_i                 : in  std_logic;  -- dahlia_fpga_awready_axi_s2_o
    fabric_fpga_bid_axi_s2_i1                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i2                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i3                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i4                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i5                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i6                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i7                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i8                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i9                    : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i10                   : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i11                   : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bid_axi_s2_i12                   : in  std_logic;  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bresp_axi_s2_i1                  : in  std_logic;  -- dahlia_fpga_bresp_axi_s2_o
    fabric_fpga_bresp_axi_s2_i2                  : in  std_logic;  -- dahlia_fpga_bresp_axi_s2_o
    fabric_fpga_bvalid_axi_s2_i                  : in  std_logic;  -- dahlia_fpga_bvalid_axi_s2_o
    fabric_fpga_rdata_axi_s2_i1                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i2                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i3                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i4                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i5                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i6                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i7                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i8                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i9                  : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i10                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i11                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i12                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i13                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i14                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i15                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i16                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i17                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i18                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i19                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i20                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i21                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i22                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i23                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i24                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i25                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i26                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i27                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i28                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i29                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i30                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i31                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i32                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i33                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i34                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i35                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i36                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i37                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i38                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i39                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i40                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i41                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i42                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i43                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i44                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i45                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i46                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i47                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i48                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i49                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i50                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i51                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i52                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i53                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i54                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i55                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i56                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i57                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i58                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i59                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i60                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i61                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i62                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i63                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i64                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i65                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i66                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i67                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i68                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i69                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i70                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i71                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i72                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i73                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i74                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i75                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i76                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i77                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i78                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i79                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i80                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i81                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i82                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i83                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i84                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i85                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i86                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i87                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i88                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i89                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i90                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i91                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i92                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i93                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i94                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i95                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i96                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i97                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i98                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i99                 : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i100                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i101                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i102                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i103                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i104                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i105                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i106                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i107                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i108                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i109                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i110                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i111                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i112                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i113                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i114                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i115                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i116                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i117                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i118                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i119                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i120                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i121                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i122                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i123                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i124                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i125                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i126                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i127                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rdata_axi_s2_i128                : in  std_logic;  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rid_axi_s2_i1                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i2                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i3                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i4                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i5                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i6                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i7                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i8                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i9                    : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i10                   : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i11                   : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rid_axi_s2_i12                   : in  std_logic;  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rlast_axi_s2_i                   : in  std_logic;  -- dahlia_fpga_rlast_axi_s2_o
    fabric_fpga_rresp_axi_s2_i1                  : in  std_logic;  -- dahlia_fpga_rresp_axi_s2_o
    fabric_fpga_rresp_axi_s2_i2                  : in  std_logic;  -- dahlia_fpga_rresp_axi_s2_o
    fabric_fpga_rvalid_axi_s2_i                  : in  std_logic;  -- dahlia_fpga_rvalid_axi_s2_o
    fabric_fpga_wready_axi_s2_i                  : in  std_logic;  -- dahlia_fpga_wready_axi_s2_o
    fabric_fpga_arready_axi_m1_o                 : out std_logic;  -- dahlia_fpga_arready_axi_m1_i
    fabric_fpga_awready_axi_m1_o                 : out std_logic;  -- dahlia_fpga_awready_axi_m1_i
    fabric_fpga_bid_axi_m1_o1                    : out std_logic;  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bid_axi_m1_o2                    : out std_logic;  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bid_axi_m1_o3                    : out std_logic;  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bid_axi_m1_o4                    : out std_logic;  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bid_axi_m1_o5                    : out std_logic;  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bresp_axi_m1_o1                  : out std_logic;  -- dahlia_fpga_bresp_axi_m1_i
    fabric_fpga_bresp_axi_m1_o2                  : out std_logic;  -- dahlia_fpga_bresp_axi_m1_i
    fabric_fpga_bvalid_axi_m1_o                  : out std_logic;  -- dahlia_fpga_bvalid_axi_m1_i
    fabric_fpga_dma_ack_m1_o1                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_ack_m1_o2                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_ack_m1_o3                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_ack_m1_o4                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_ack_m1_o5                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_ack_m1_o6                    : out std_logic;  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_finish_m1_o1                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_dma_finish_m1_o2                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_dma_finish_m1_o3                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_dma_finish_m1_o4                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_dma_finish_m1_o5                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_dma_finish_m1_o6                 : out std_logic;  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_rdata_axi_m1_o1                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o2                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o3                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o4                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o5                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o6                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o7                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o8                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o9                  : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o10                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o11                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o12                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o13                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o14                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o15                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o16                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o17                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o18                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o19                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o20                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o21                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o22                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o23                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o24                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o25                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o26                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o27                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o28                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o29                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o30                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o31                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o32                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o33                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o34                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o35                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o36                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o37                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o38                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o39                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o40                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o41                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o42                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o43                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o44                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o45                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o46                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o47                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o48                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o49                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o50                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o51                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o52                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o53                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o54                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o55                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o56                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o57                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o58                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o59                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o60                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o61                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o62                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o63                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o64                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o65                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o66                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o67                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o68                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o69                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o70                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o71                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o72                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o73                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o74                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o75                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o76                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o77                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o78                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o79                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o80                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o81                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o82                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o83                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o84                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o85                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o86                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o87                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o88                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o89                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o90                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o91                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o92                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o93                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o94                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o95                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o96                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o97                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o98                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o99                 : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o100                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o101                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o102                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o103                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o104                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o105                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o106                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o107                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o108                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o109                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o110                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o111                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o112                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o113                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o114                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o115                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o116                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o117                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o118                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o119                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o120                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o121                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o122                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o123                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o124                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o125                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o126                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o127                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rdata_axi_m1_o128                : out std_logic;  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rid_axi_m1_o1                    : out std_logic;  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rid_axi_m1_o2                    : out std_logic;  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rid_axi_m1_o3                    : out std_logic;  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rid_axi_m1_o4                    : out std_logic;  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rid_axi_m1_o5                    : out std_logic;  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rlast_axi_m1_o                   : out std_logic;  -- dahlia_fpga_rlast_axi_m1_i
    fabric_fpga_rresp_axi_m1_o1                  : out std_logic;  -- dahlia_fpga_rresp_axi_m1_i
    fabric_fpga_rresp_axi_m1_o2                  : out std_logic;  -- dahlia_fpga_rresp_axi_m1_i
    fabric_fpga_rvalid_axi_m1_o                  : out std_logic;  -- dahlia_fpga_rvalid_axi_m1_i
    fabric_fpga_wready_axi_m1_o                  : out std_logic;  -- dahlia_fpga_wready_axi_m1_i
    fabric_fpga_araddr_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i4                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i5                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i6                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i7                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i8                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i9                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i10                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i11                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i12                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i13                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i14                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i15                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i16                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i17                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i18                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i19                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i20                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i21                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i22                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i23                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i24                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i25                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i26                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i27                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i28                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i29                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i30                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i31                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i32                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i33                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i34                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i35                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i36                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i37                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i38                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i39                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_araddr_axi_m1_i40                : in  std_logic;  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_arburst_axi_m1_i1                : in  std_logic;  -- dahlia_fpga_arburst_axi_m1_o
    fabric_fpga_arburst_axi_m1_i2                : in  std_logic;  -- dahlia_fpga_arburst_axi_m1_o
    fabric_fpga_arcache_axi_m1_i1                : in  std_logic;  -- dahlia_fpga_arcache_axi_m1_o
    fabric_fpga_arcache_axi_m1_i2                : in  std_logic;  -- dahlia_fpga_arcache_axi_m1_o
    fabric_fpga_arcache_axi_m1_i3                : in  std_logic;  -- dahlia_fpga_arcache_axi_m1_o
    fabric_fpga_arcache_axi_m1_i4                : in  std_logic;  -- dahlia_fpga_arcache_axi_m1_o
    fabric_fpga_arid_axi_m1_i1                   : in  std_logic;  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arid_axi_m1_i2                   : in  std_logic;  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arid_axi_m1_i3                   : in  std_logic;  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arid_axi_m1_i4                   : in  std_logic;  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arid_axi_m1_i5                   : in  std_logic;  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arlen_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i5                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i6                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i7                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlen_axi_m1_i8                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlock_axi_m1_i                  : in  std_logic;  -- dahlia_fpga_arlock_axi_m1_o
    fabric_fpga_arprot_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m1_o
    fabric_fpga_arprot_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m1_o
    fabric_fpga_arprot_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m1_o
    fabric_fpga_arqos_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m1_o
    fabric_fpga_arqos_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m1_o
    fabric_fpga_arqos_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m1_o
    fabric_fpga_arqos_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m1_o
    fabric_fpga_arsize_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m1_o
    fabric_fpga_arsize_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m1_o
    fabric_fpga_arsize_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m1_o
    fabric_fpga_arvalid_axi_m1_i                 : in  std_logic;  -- dahlia_fpga_arvalid_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i4                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i5                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i6                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i7                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i8                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i9                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i10                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i11                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i12                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i13                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i14                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i15                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i16                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i17                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i18                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i19                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i20                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i21                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i22                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i23                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i24                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i25                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i26                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i27                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i28                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i29                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i30                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i31                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i32                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i33                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i34                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i35                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i36                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i37                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i38                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i39                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i40                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awburst_axi_m1_i1                : in  std_logic;  -- dahlia_fpga_awburst_axi_m1_o
    fabric_fpga_awburst_axi_m1_i2                : in  std_logic;  -- dahlia_fpga_awburst_axi_m1_o
    fabric_fpga_awcache_axi_m1_i1                : in  std_logic;  -- dahlia_fpga_awcache_axi_m1_o
    fabric_fpga_awcache_axi_m1_i2                : in  std_logic;  -- dahlia_fpga_awcache_axi_m1_o
    fabric_fpga_awcache_axi_m1_i3                : in  std_logic;  -- dahlia_fpga_awcache_axi_m1_o
    fabric_fpga_awcache_axi_m1_i4                : in  std_logic;  -- dahlia_fpga_awcache_axi_m1_o
    fabric_fpga_awid_axi_m1_i1                   : in  std_logic;  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awid_axi_m1_i2                   : in  std_logic;  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awid_axi_m1_i3                   : in  std_logic;  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awid_axi_m1_i4                   : in  std_logic;  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awid_axi_m1_i5                   : in  std_logic;  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awlen_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i5                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i6                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i7                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlen_axi_m1_i8                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlock_axi_m1_i                  : in  std_logic;  -- dahlia_fpga_awlock_axi_m1_o
    fabric_fpga_awprot_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m1_o
    fabric_fpga_awprot_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m1_o
    fabric_fpga_awprot_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m1_o
    fabric_fpga_awqos_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m1_o
    fabric_fpga_awqos_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m1_o
    fabric_fpga_awqos_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m1_o
    fabric_fpga_awqos_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m1_o
    fabric_fpga_awsize_axi_m1_i1                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m1_o
    fabric_fpga_awsize_axi_m1_i2                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m1_o
    fabric_fpga_awsize_axi_m1_i3                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m1_o
    fabric_fpga_awvalid_axi_m1_i                 : in  std_logic;  -- dahlia_fpga_awvalid_axi_m1_o
    fabric_fpga_bready_axi_m1_i                  : in  std_logic;  -- dahlia_fpga_bready_axi_m1_o
    fabric_fpga_dma_last_m1_i1                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_last_m1_i2                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_last_m1_i3                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_last_m1_i4                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_last_m1_i5                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_last_m1_i6                   : in  std_logic;  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_req_m1_i1                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_req_m1_i2                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_req_m1_i3                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_req_m1_i4                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_req_m1_i5                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_req_m1_i6                    : in  std_logic;  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_single_m1_i1                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_dma_single_m1_i2                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_dma_single_m1_i3                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_dma_single_m1_i4                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_dma_single_m1_i5                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_dma_single_m1_i6                 : in  std_logic;  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_rready_axi_m1_i                  : in  std_logic;  -- dahlia_fpga_rready_axi_m1_o
    fabric_fpga_wdata_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i5                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i6                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i7                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i8                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i9                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i10                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i11                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i12                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i13                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i14                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i15                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i16                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i17                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i18                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i19                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i20                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i21                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i22                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i23                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i24                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i25                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i26                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i27                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i28                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i29                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i30                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i31                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i32                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i33                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i34                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i35                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i36                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i37                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i38                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i39                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i40                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i41                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i42                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i43                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i44                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i45                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i46                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i47                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i48                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i49                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i50                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i51                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i52                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i53                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i54                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i55                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i56                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i57                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i58                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i59                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i60                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i61                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i62                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i63                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i64                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i65                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i66                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i67                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i68                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i69                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i70                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i71                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i72                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i73                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i74                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i75                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i76                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i77                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i78                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i79                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i80                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i81                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i82                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i83                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i84                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i85                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i86                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i87                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i88                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i89                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i90                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i91                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i92                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i93                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i94                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i95                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i96                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i97                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i98                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i99                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i100                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i101                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i102                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i103                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i104                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i105                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i106                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i107                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i108                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i109                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i110                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i111                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i112                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i113                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i114                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i115                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i116                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i117                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i118                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i119                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i120                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i121                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i122                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i123                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i124                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i125                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i126                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i127                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wdata_axi_m1_i128                : in  std_logic;  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wlast_axi_m1_i                   : in  std_logic;  -- dahlia_fpga_wlast_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i1                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i2                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i3                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i4                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i5                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i6                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i7                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i8                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i9                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i10                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i11                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i12                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i13                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i14                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i15                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i16                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wvalid_axi_m1_i                  : in  std_logic;  -- dahlia_fpga_wvalid_axi_m1_o
    fabric_fpga_arready_axi_m2_o                 : out std_logic;  -- dahlia_fpga_arready_axi_m2_i
    fabric_fpga_awready_axi_m2_o                 : out std_logic;  -- dahlia_fpga_awready_axi_m2_i
    fabric_fpga_bid_axi_m2_o1                    : out std_logic;  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bid_axi_m2_o2                    : out std_logic;  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bid_axi_m2_o3                    : out std_logic;  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bid_axi_m2_o4                    : out std_logic;  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bid_axi_m2_o5                    : out std_logic;  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bresp_axi_m2_o1                  : out std_logic;  -- dahlia_fpga_bresp_axi_m2_i
    fabric_fpga_bresp_axi_m2_o2                  : out std_logic;  -- dahlia_fpga_bresp_axi_m2_i
    fabric_fpga_bvalid_axi_m2_o                  : out std_logic;  -- dahlia_fpga_bvalid_axi_m2_i
    fabric_fpga_dma_ack_m2_o1                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_ack_m2_o2                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_ack_m2_o3                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_ack_m2_o4                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_ack_m2_o5                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_ack_m2_o6                    : out std_logic;  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_finish_m2_o1                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_dma_finish_m2_o2                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_dma_finish_m2_o3                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_dma_finish_m2_o4                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_dma_finish_m2_o5                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_dma_finish_m2_o6                 : out std_logic;  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_rdata_axi_m2_o1                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o2                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o3                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o4                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o5                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o6                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o7                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o8                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o9                  : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o10                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o11                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o12                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o13                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o14                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o15                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o16                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o17                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o18                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o19                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o20                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o21                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o22                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o23                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o24                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o25                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o26                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o27                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o28                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o29                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o30                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o31                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o32                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o33                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o34                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o35                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o36                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o37                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o38                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o39                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o40                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o41                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o42                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o43                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o44                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o45                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o46                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o47                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o48                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o49                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o50                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o51                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o52                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o53                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o54                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o55                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o56                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o57                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o58                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o59                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o60                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o61                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o62                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o63                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o64                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o65                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o66                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o67                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o68                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o69                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o70                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o71                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o72                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o73                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o74                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o75                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o76                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o77                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o78                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o79                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o80                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o81                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o82                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o83                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o84                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o85                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o86                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o87                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o88                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o89                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o90                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o91                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o92                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o93                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o94                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o95                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o96                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o97                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o98                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o99                 : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o100                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o101                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o102                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o103                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o104                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o105                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o106                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o107                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o108                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o109                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o110                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o111                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o112                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o113                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o114                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o115                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o116                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o117                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o118                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o119                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o120                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o121                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o122                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o123                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o124                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o125                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o126                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o127                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rdata_axi_m2_o128                : out std_logic;  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rid_axi_m2_o1                    : out std_logic;  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rid_axi_m2_o2                    : out std_logic;  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rid_axi_m2_o3                    : out std_logic;  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rid_axi_m2_o4                    : out std_logic;  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rid_axi_m2_o5                    : out std_logic;  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rlast_axi_m2_o                   : out std_logic;  -- dahlia_fpga_rlast_axi_m2_i
    fabric_fpga_rresp_axi_m2_o1                  : out std_logic;  -- dahlia_fpga_rresp_axi_m2_i
    fabric_fpga_rresp_axi_m2_o2                  : out std_logic;  -- dahlia_fpga_rresp_axi_m2_i
    fabric_fpga_rvalid_axi_m2_o                  : out std_logic;  -- dahlia_fpga_rvalid_axi_m2_i
    fabric_fpga_wready_axi_m2_o                  : out std_logic;  -- dahlia_fpga_wready_axi_m2_i
    fabric_fpga_araddr_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i4                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i5                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i6                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i7                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i8                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i9                 : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i10                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i11                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i12                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i13                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i14                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i15                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i16                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i17                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i18                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i19                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i20                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i21                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i22                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i23                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i24                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i25                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i26                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i27                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i28                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i29                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i30                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i31                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i32                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i33                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i34                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i35                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i36                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i37                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i38                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i39                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_araddr_axi_m2_i40                : in  std_logic;  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_arburst_axi_m2_i1                : in  std_logic;  -- dahlia_fpga_arburst_axi_m2_o
    fabric_fpga_arburst_axi_m2_i2                : in  std_logic;  -- dahlia_fpga_arburst_axi_m2_o
    fabric_fpga_arcache_axi_m2_i1                : in  std_logic;  -- dahlia_fpga_arcache_axi_m2_o
    fabric_fpga_arcache_axi_m2_i2                : in  std_logic;  -- dahlia_fpga_arcache_axi_m2_o
    fabric_fpga_arcache_axi_m2_i3                : in  std_logic;  -- dahlia_fpga_arcache_axi_m2_o
    fabric_fpga_arcache_axi_m2_i4                : in  std_logic;  -- dahlia_fpga_arcache_axi_m2_o
    fabric_fpga_arid_axi_m2_i1                   : in  std_logic;  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arid_axi_m2_i2                   : in  std_logic;  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arid_axi_m2_i3                   : in  std_logic;  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arid_axi_m2_i4                   : in  std_logic;  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arid_axi_m2_i5                   : in  std_logic;  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arlen_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i5                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i6                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i7                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlen_axi_m2_i8                  : in  std_logic;  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlock_axi_m2_i                  : in  std_logic;  -- dahlia_fpga_arlock_axi_m2_o
    fabric_fpga_arprot_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m2_o
    fabric_fpga_arprot_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m2_o
    fabric_fpga_arprot_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_arprot_axi_m2_o
    fabric_fpga_arqos_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m2_o
    fabric_fpga_arqos_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m2_o
    fabric_fpga_arqos_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m2_o
    fabric_fpga_arqos_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_arqos_axi_m2_o
    fabric_fpga_arsize_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m2_o
    fabric_fpga_arsize_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m2_o
    fabric_fpga_arsize_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_arsize_axi_m2_o
    fabric_fpga_arvalid_axi_m2_i                 : in  std_logic;  -- dahlia_fpga_arvalid_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i4                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i5                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i6                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i7                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i8                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i9                 : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i10                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i11                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i12                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i13                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i14                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i15                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i16                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i17                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i18                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i19                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i20                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i21                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i22                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i23                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i24                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i25                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i26                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i27                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i28                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i29                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i30                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i31                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i32                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i33                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i34                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i35                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i36                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i37                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i38                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i39                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i40                : in  std_logic;  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awburst_axi_m2_i1                : in  std_logic;  -- dahlia_fpga_awburst_axi_m2_o
    fabric_fpga_awburst_axi_m2_i2                : in  std_logic;  -- dahlia_fpga_awburst_axi_m2_o
    fabric_fpga_awcache_axi_m2_i1                : in  std_logic;  -- dahlia_fpga_awcache_axi_m2_o
    fabric_fpga_awcache_axi_m2_i2                : in  std_logic;  -- dahlia_fpga_awcache_axi_m2_o
    fabric_fpga_awcache_axi_m2_i3                : in  std_logic;  -- dahlia_fpga_awcache_axi_m2_o
    fabric_fpga_awcache_axi_m2_i4                : in  std_logic;  -- dahlia_fpga_awcache_axi_m2_o
    fabric_fpga_awid_axi_m2_i1                   : in  std_logic;  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awid_axi_m2_i2                   : in  std_logic;  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awid_axi_m2_i3                   : in  std_logic;  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awid_axi_m2_i4                   : in  std_logic;  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awid_axi_m2_i5                   : in  std_logic;  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awlen_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i5                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i6                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i7                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlen_axi_m2_i8                  : in  std_logic;  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlock_axi_m2_i                  : in  std_logic;  -- dahlia_fpga_awlock_axi_m2_o
    fabric_fpga_awprot_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m2_o
    fabric_fpga_awprot_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m2_o
    fabric_fpga_awprot_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_awprot_axi_m2_o
    fabric_fpga_awqos_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m2_o
    fabric_fpga_awqos_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m2_o
    fabric_fpga_awqos_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m2_o
    fabric_fpga_awqos_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_awqos_axi_m2_o
    fabric_fpga_awsize_axi_m2_i1                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m2_o
    fabric_fpga_awsize_axi_m2_i2                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m2_o
    fabric_fpga_awsize_axi_m2_i3                 : in  std_logic;  -- dahlia_fpga_awsize_axi_m2_o
    fabric_fpga_awvalid_axi_m2_i                 : in  std_logic;  -- dahlia_fpga_awvalid_axi_m2_o
    fabric_fpga_bready_axi_m2_i                  : in  std_logic;  -- dahlia_fpga_bready_axi_m2_o
    fabric_fpga_dma_last_m2_i1                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_last_m2_i2                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_last_m2_i3                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_last_m2_i4                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_last_m2_i5                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_last_m2_i6                   : in  std_logic;  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_req_m2_i1                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_req_m2_i2                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_req_m2_i3                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_req_m2_i4                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_req_m2_i5                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_req_m2_i6                    : in  std_logic;  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_single_m2_i1                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_dma_single_m2_i2                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_dma_single_m2_i3                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_dma_single_m2_i4                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_dma_single_m2_i5                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_dma_single_m2_i6                 : in  std_logic;  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_rready_axi_m2_i                  : in  std_logic;  -- dahlia_fpga_rready_axi_m2_o
    fabric_fpga_wdata_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i5                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i6                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i7                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i8                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i9                  : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i10                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i11                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i12                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i13                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i14                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i15                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i16                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i17                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i18                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i19                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i20                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i21                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i22                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i23                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i24                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i25                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i26                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i27                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i28                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i29                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i30                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i31                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i32                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i33                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i34                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i35                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i36                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i37                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i38                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i39                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i40                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i41                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i42                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i43                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i44                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i45                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i46                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i47                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i48                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i49                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i50                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i51                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i52                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i53                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i54                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i55                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i56                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i57                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i58                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i59                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i60                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i61                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i62                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i63                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i64                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i65                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i66                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i67                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i68                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i69                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i70                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i71                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i72                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i73                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i74                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i75                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i76                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i77                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i78                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i79                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i80                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i81                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i82                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i83                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i84                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i85                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i86                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i87                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i88                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i89                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i90                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i91                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i92                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i93                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i94                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i95                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i96                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i97                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i98                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i99                 : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i100                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i101                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i102                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i103                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i104                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i105                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i106                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i107                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i108                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i109                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i110                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i111                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i112                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i113                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i114                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i115                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i116                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i117                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i118                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i119                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i120                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i121                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i122                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i123                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i124                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i125                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i126                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i127                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wdata_axi_m2_i128                : in  std_logic;  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wlast_axi_m2_i                   : in  std_logic;  -- dahlia_fpga_wlast_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i1                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i2                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i3                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i4                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i5                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i6                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i7                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i8                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i9                  : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i10                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i11                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i12                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i13                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i14                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i15                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i16                 : in  std_logic;  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wvalid_axi_m2_i                  : in  std_logic;  -- dahlia_fpga_wvalid_axi_m2_o
    fabric_fpga_ddr0_arready_o                   : out std_logic;  -- dahlia_fpga_ddr0_arready_i
    fabric_fpga_ddr0_awready_o                   : out std_logic;  -- dahlia_fpga_ddr0_awready_i
    fabric_fpga_ddr0_bid_o1                      : out std_logic;  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bid_o2                      : out std_logic;  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bid_o3                      : out std_logic;  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bid_o4                      : out std_logic;  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bid_o5                      : out std_logic;  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bresp_o1                    : out std_logic;  -- dahlia_fpga_ddr0_bresp_i
    fabric_fpga_ddr0_bresp_o2                    : out std_logic;  -- dahlia_fpga_ddr0_bresp_i
    fabric_fpga_ddr0_bvalid_o                    : out std_logic;  -- dahlia_fpga_ddr0_bvalid_i
    fabric_fpga_ddr0_rdata_o1                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o2                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o3                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o4                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o5                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o6                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o7                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o8                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o9                    : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o10                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o11                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o12                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o13                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o14                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o15                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o16                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o17                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o18                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o19                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o20                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o21                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o22                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o23                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o24                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o25                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o26                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o27                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o28                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o29                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o30                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o31                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o32                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o33                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o34                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o35                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o36                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o37                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o38                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o39                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o40                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o41                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o42                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o43                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o44                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o45                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o46                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o47                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o48                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o49                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o50                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o51                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o52                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o53                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o54                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o55                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o56                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o57                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o58                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o59                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o60                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o61                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o62                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o63                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o64                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o65                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o66                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o67                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o68                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o69                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o70                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o71                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o72                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o73                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o74                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o75                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o76                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o77                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o78                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o79                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o80                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o81                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o82                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o83                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o84                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o85                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o86                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o87                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o88                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o89                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o90                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o91                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o92                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o93                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o94                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o95                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o96                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o97                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o98                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o99                   : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o100                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o101                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o102                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o103                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o104                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o105                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o106                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o107                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o108                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o109                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o110                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o111                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o112                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o113                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o114                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o115                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o116                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o117                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o118                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o119                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o120                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o121                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o122                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o123                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o124                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o125                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o126                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o127                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rdata_o128                  : out std_logic;  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rid_o1                      : out std_logic;  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rid_o2                      : out std_logic;  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rid_o3                      : out std_logic;  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rid_o4                      : out std_logic;  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rid_o5                      : out std_logic;  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rlast_o                     : out std_logic;  -- dahlia_fpga_ddr0_rlast_i
    fabric_fpga_ddr0_rresp_o1                    : out std_logic;  -- dahlia_fpga_ddr0_rresp_i
    fabric_fpga_ddr0_rresp_o2                    : out std_logic;  -- dahlia_fpga_ddr0_rresp_i
    fabric_fpga_ddr0_rvalid_o                    : out std_logic;  -- dahlia_fpga_ddr0_rvalid_i
    fabric_fpga_ddr0_wready_o                    : out std_logic;  -- dahlia_fpga_ddr0_wready_i
    fabric_fpga_ddr0_araddr_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i4                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i5                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i6                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i7                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i8                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i9                   : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i10                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i11                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i12                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i13                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i14                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i15                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i16                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i17                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i18                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i19                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i20                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i21                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i22                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i23                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i24                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i25                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i26                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i27                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i28                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i29                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i30                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i31                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i32                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i33                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i34                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i35                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i36                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i37                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i38                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i39                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_araddr_i40                  : in  std_logic;  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_arburst_i1                  : in  std_logic;  -- dahlia_fpga_ddr0_arburst_o
    fabric_fpga_ddr0_arburst_i2                  : in  std_logic;  -- dahlia_fpga_ddr0_arburst_o
    fabric_fpga_ddr0_arcache_i1                  : in  std_logic;  -- dahlia_fpga_ddr0_arcache_o
    fabric_fpga_ddr0_arcache_i2                  : in  std_logic;  -- dahlia_fpga_ddr0_arcache_o
    fabric_fpga_ddr0_arcache_i3                  : in  std_logic;  -- dahlia_fpga_ddr0_arcache_o
    fabric_fpga_ddr0_arcache_i4                  : in  std_logic;  -- dahlia_fpga_ddr0_arcache_o
    fabric_fpga_ddr0_arid_i1                     : in  std_logic;  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arid_i2                     : in  std_logic;  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arid_i3                     : in  std_logic;  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arid_i4                     : in  std_logic;  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arid_i5                     : in  std_logic;  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arlen_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i5                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i6                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i7                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlen_i8                    : in  std_logic;  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlock_i                    : in  std_logic;  -- dahlia_fpga_ddr0_arlock_o
    fabric_fpga_ddr0_arprot_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_arprot_o
    fabric_fpga_ddr0_arprot_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_arprot_o
    fabric_fpga_ddr0_arprot_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_arprot_o
    fabric_fpga_ddr0_arqos_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_arqos_o
    fabric_fpga_ddr0_arqos_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_arqos_o
    fabric_fpga_ddr0_arqos_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_arqos_o
    fabric_fpga_ddr0_arqos_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_arqos_o
    fabric_fpga_ddr0_arsize_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_arsize_o
    fabric_fpga_ddr0_arsize_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_arsize_o
    fabric_fpga_ddr0_arsize_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_arsize_o
    fabric_fpga_ddr0_arvalid_i                   : in  std_logic;  -- dahlia_fpga_ddr0_arvalid_o
    fabric_fpga_ddr0_awaddr_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i4                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i5                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i6                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i7                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i8                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i9                   : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i10                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i11                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i12                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i13                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i14                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i15                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i16                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i17                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i18                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i19                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i20                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i21                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i22                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i23                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i24                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i25                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i26                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i27                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i28                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i29                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i30                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i31                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i32                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i33                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i34                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i35                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i36                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i37                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i38                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i39                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awaddr_i40                  : in  std_logic;  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awburst_i1                  : in  std_logic;  -- dahlia_fpga_ddr0_awburst_o
    fabric_fpga_ddr0_awburst_i2                  : in  std_logic;  -- dahlia_fpga_ddr0_awburst_o
    fabric_fpga_ddr0_awcache_i1                  : in  std_logic;  -- dahlia_fpga_ddr0_awcache_o
    fabric_fpga_ddr0_awcache_i2                  : in  std_logic;  -- dahlia_fpga_ddr0_awcache_o
    fabric_fpga_ddr0_awcache_i3                  : in  std_logic;  -- dahlia_fpga_ddr0_awcache_o
    fabric_fpga_ddr0_awcache_i4                  : in  std_logic;  -- dahlia_fpga_ddr0_awcache_o
    fabric_fpga_ddr0_awid_i1                     : in  std_logic;  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awid_i2                     : in  std_logic;  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awid_i3                     : in  std_logic;  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awid_i4                     : in  std_logic;  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awid_i5                     : in  std_logic;  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awlen_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i5                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i6                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i7                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlen_i8                    : in  std_logic;  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlock_i                    : in  std_logic;  -- dahlia_fpga_ddr0_awlock_o
    fabric_fpga_ddr0_awprot_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_awprot_o
    fabric_fpga_ddr0_awprot_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_awprot_o
    fabric_fpga_ddr0_awprot_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_awprot_o
    fabric_fpga_ddr0_awqos_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_awqos_o
    fabric_fpga_ddr0_awqos_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_awqos_o
    fabric_fpga_ddr0_awqos_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_awqos_o
    fabric_fpga_ddr0_awqos_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_awqos_o
    fabric_fpga_ddr0_awsize_i1                   : in  std_logic;  -- dahlia_fpga_ddr0_awsize_o
    fabric_fpga_ddr0_awsize_i2                   : in  std_logic;  -- dahlia_fpga_ddr0_awsize_o
    fabric_fpga_ddr0_awsize_i3                   : in  std_logic;  -- dahlia_fpga_ddr0_awsize_o
    fabric_fpga_ddr0_awvalid_i                   : in  std_logic;  -- dahlia_fpga_ddr0_awvalid_o
    fabric_fpga_ddr0_bready_i                    : in  std_logic;  -- dahlia_fpga_ddr0_bready_o
    fabric_fpga_ddr0_rready_i                    : in  std_logic;  -- dahlia_fpga_ddr0_rready_o
    fabric_fpga_ddr0_wdata_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i5                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i6                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i7                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i8                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i9                    : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i10                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i11                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i12                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i13                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i14                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i15                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i16                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i17                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i18                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i19                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i20                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i21                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i22                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i23                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i24                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i25                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i26                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i27                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i28                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i29                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i30                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i31                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i32                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i33                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i34                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i35                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i36                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i37                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i38                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i39                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i40                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i41                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i42                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i43                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i44                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i45                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i46                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i47                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i48                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i49                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i50                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i51                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i52                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i53                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i54                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i55                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i56                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i57                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i58                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i59                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i60                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i61                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i62                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i63                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i64                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i65                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i66                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i67                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i68                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i69                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i70                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i71                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i72                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i73                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i74                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i75                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i76                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i77                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i78                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i79                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i80                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i81                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i82                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i83                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i84                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i85                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i86                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i87                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i88                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i89                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i90                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i91                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i92                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i93                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i94                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i95                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i96                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i97                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i98                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i99                   : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i100                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i101                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i102                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i103                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i104                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i105                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i106                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i107                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i108                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i109                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i110                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i111                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i112                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i113                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i114                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i115                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i116                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i117                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i118                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i119                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i120                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i121                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i122                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i123                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i124                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i125                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i126                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i127                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wdata_i128                  : in  std_logic;  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wlast_i                     : in  std_logic;  -- dahlia_fpga_ddr0_wlast_o
    fabric_fpga_ddr0_wstrb_i1                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i2                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i3                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i4                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i5                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i6                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i7                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i8                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i9                    : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i10                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i11                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i12                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i13                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i14                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i15                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wstrb_i16                   : in  std_logic;  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wvalid_i                    : in  std_logic;  -- dahlia_fpga_ddr0_wvalid_o
    fabric_fpga_paddr_apb_o1                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o2                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o3                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o4                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o5                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o6                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o7                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o8                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o9                     : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o10                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o11                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o12                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o13                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o14                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o15                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o16                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o17                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o18                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o19                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o20                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o21                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o22                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o23                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o24                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o25                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o26                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o27                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o28                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o29                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o30                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o31                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_paddr_apb_o32                    : out std_logic;  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_penable_apb_o                    : out std_logic;  -- dahlia_fpga_penable_apb_i
    fabric_fpga_psel_apb_o                       : out std_logic;  -- dahlia_fpga_psel_apb_i
    fabric_fpga_pwdata_apb_o1                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o2                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o3                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o4                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o5                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o6                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o7                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o8                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o9                    : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o10                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o11                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o12                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o13                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o14                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o15                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o16                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o17                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o18                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o19                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o20                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o21                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o22                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o23                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o24                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o25                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o26                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o27                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o28                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o29                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o30                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o31                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwdata_apb_o32                   : out std_logic;  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwrite_apb_o                     : out std_logic;  -- dahlia_fpga_pwrite_apb_i
    fabric_fpga_prdata_apb_i1                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i2                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i3                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i4                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i5                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i6                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i7                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i8                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i9                    : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i10                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i11                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i12                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i13                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i14                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i15                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i16                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i17                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i18                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i19                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i20                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i21                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i22                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i23                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i24                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i25                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i26                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i27                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i28                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i29                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i30                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i31                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_prdata_apb_i32                   : in  std_logic;  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_pready_apb_i                     : in  std_logic;  -- dahlia_fpga_pready_apb_o
    fabric_fpga_pslverr_apb_i                    : in  std_logic;  -- dahlia_fpga_pslverr_apb_o
    fabric_llpp0_araddr_s_o1                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o2                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o3                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o4                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o5                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o6                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o7                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o8                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o9                     : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o10                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o11                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o12                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o13                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o14                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o15                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o16                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o17                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o18                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o19                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o20                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o21                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o22                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o23                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o24                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o25                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o26                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o27                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o28                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o29                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o30                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o31                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_araddr_s_o32                    : out std_logic;  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_arburst_s_o1                    : out std_logic;  -- dahlia_llpp0_arburst_s_i
    fabric_llpp0_arburst_s_o2                    : out std_logic;  -- dahlia_llpp0_arburst_s_i
    fabric_llpp0_arcache_s_o1                    : out std_logic;  -- dahlia_llpp0_arcache_s_i
    fabric_llpp0_arcache_s_o2                    : out std_logic;  -- dahlia_llpp0_arcache_s_i
    fabric_llpp0_arcache_s_o3                    : out std_logic;  -- dahlia_llpp0_arcache_s_i
    fabric_llpp0_arcache_s_o4                    : out std_logic;  -- dahlia_llpp0_arcache_s_i
    fabric_llpp0_arid_s_o1                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o2                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o3                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o4                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o5                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o6                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o7                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o8                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o9                       : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o10                      : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o11                      : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arid_s_o12                      : out std_logic;  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arlen_s_o1                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o2                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o3                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o4                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o5                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o6                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o7                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlen_s_o8                      : out std_logic;  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlock_s_o                      : out std_logic;  -- dahlia_llpp0_arlock_s_i
    fabric_llpp0_arprot_s_o1                     : out std_logic;  -- dahlia_llpp0_arprot_s_i
    fabric_llpp0_arprot_s_o2                     : out std_logic;  -- dahlia_llpp0_arprot_s_i
    fabric_llpp0_arprot_s_o3                     : out std_logic;  -- dahlia_llpp0_arprot_s_i
    fabric_llpp0_arqos_s_o1                      : out std_logic;  -- dahlia_llpp0_arqos_s_i
    fabric_llpp0_arqos_s_o2                      : out std_logic;  -- dahlia_llpp0_arqos_s_i
    fabric_llpp0_arqos_s_o3                      : out std_logic;  -- dahlia_llpp0_arqos_s_i
    fabric_llpp0_arqos_s_o4                      : out std_logic;  -- dahlia_llpp0_arqos_s_i
    fabric_llpp0_arsize_s_o1                     : out std_logic;  -- dahlia_llpp0_arsize_s_i
    fabric_llpp0_arsize_s_o2                     : out std_logic;  -- dahlia_llpp0_arsize_s_i
    fabric_llpp0_arsize_s_o3                     : out std_logic;  -- dahlia_llpp0_arsize_s_i
    fabric_llpp0_arvalid_s_o                     : out std_logic;  -- dahlia_llpp0_arvalid_s_i
    fabric_llpp0_awaddr_s_o1                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o2                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o3                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o4                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o5                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o6                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o7                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o8                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o9                     : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o10                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o11                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o12                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o13                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o14                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o15                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o16                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o17                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o18                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o19                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o20                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o21                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o22                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o23                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o24                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o25                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o26                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o27                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o28                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o29                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o30                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o31                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awaddr_s_o32                    : out std_logic;  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awburst_s_o1                    : out std_logic;  -- dahlia_llpp0_awburst_s_i
    fabric_llpp0_awburst_s_o2                    : out std_logic;  -- dahlia_llpp0_awburst_s_i
    fabric_llpp0_awcache_s_o1                    : out std_logic;  -- dahlia_llpp0_awcache_s_i
    fabric_llpp0_awcache_s_o2                    : out std_logic;  -- dahlia_llpp0_awcache_s_i
    fabric_llpp0_awcache_s_o3                    : out std_logic;  -- dahlia_llpp0_awcache_s_i
    fabric_llpp0_awcache_s_o4                    : out std_logic;  -- dahlia_llpp0_awcache_s_i
    fabric_llpp0_awid_s_o1                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o2                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o3                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o4                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o5                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o6                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o7                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o8                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o9                       : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o10                      : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o11                      : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awid_s_o12                      : out std_logic;  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awlen_s_o1                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o2                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o3                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o4                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o5                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o6                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o7                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlen_s_o8                      : out std_logic;  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlock_s_o                      : out std_logic;  -- dahlia_llpp0_awlock_s_i
    fabric_llpp0_awprot_s_o1                     : out std_logic;  -- dahlia_llpp0_awprot_s_i
    fabric_llpp0_awprot_s_o2                     : out std_logic;  -- dahlia_llpp0_awprot_s_i
    fabric_llpp0_awprot_s_o3                     : out std_logic;  -- dahlia_llpp0_awprot_s_i
    fabric_llpp0_awqos_s_o1                      : out std_logic;  -- dahlia_llpp0_awqos_s_i
    fabric_llpp0_awqos_s_o2                      : out std_logic;  -- dahlia_llpp0_awqos_s_i
    fabric_llpp0_awqos_s_o3                      : out std_logic;  -- dahlia_llpp0_awqos_s_i
    fabric_llpp0_awqos_s_o4                      : out std_logic;  -- dahlia_llpp0_awqos_s_i
    fabric_llpp0_awsize_s_o1                     : out std_logic;  -- dahlia_llpp0_awsize_s_i
    fabric_llpp0_awsize_s_o2                     : out std_logic;  -- dahlia_llpp0_awsize_s_i
    fabric_llpp0_awsize_s_o3                     : out std_logic;  -- dahlia_llpp0_awsize_s_i
    fabric_llpp0_awvalid_s_o                     : out std_logic;  -- dahlia_llpp0_awvalid_s_i
    fabric_llpp0_bready_s_o                      : out std_logic;  -- dahlia_llpp0_bready_s_i
    fabric_llpp0_rready_s_o                      : out std_logic;  -- dahlia_llpp0_rready_s_i
    fabric_llpp0_wdata_s_o1                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o2                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o3                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o4                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o5                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o6                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o7                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o8                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o9                      : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o10                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o11                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o12                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o13                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o14                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o15                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o16                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o17                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o18                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o19                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o20                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o21                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o22                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o23                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o24                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o25                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o26                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o27                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o28                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o29                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o30                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o31                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wdata_s_o32                     : out std_logic;  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wlast_s_o                       : out std_logic;  -- dahlia_llpp0_wlast_s_i
    fabric_llpp0_wstrb_s_o1                      : out std_logic;  -- dahlia_llpp0_wstrb_s_i
    fabric_llpp0_wstrb_s_o2                      : out std_logic;  -- dahlia_llpp0_wstrb_s_i
    fabric_llpp0_wstrb_s_o3                      : out std_logic;  -- dahlia_llpp0_wstrb_s_i
    fabric_llpp0_wstrb_s_o4                      : out std_logic;  -- dahlia_llpp0_wstrb_s_i
    fabric_llpp0_wvalid_s_o                      : out std_logic;  -- dahlia_llpp0_wvalid_s_i
    fabric_llpp0_arready_s_i                     : in  std_logic;  -- dahlia_llpp0_arready_s_o
    fabric_llpp0_awready_s_i                     : in  std_logic;  -- dahlia_llpp0_awready_s_o
    fabric_llpp0_bid_s_i1                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i2                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i3                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i4                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i5                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i6                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i7                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i8                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i9                        : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i10                       : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i11                       : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bid_s_i12                       : in  std_logic;  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bresp_s_i1                      : in  std_logic;  -- dahlia_llpp0_bresp_s_o
    fabric_llpp0_bresp_s_i2                      : in  std_logic;  -- dahlia_llpp0_bresp_s_o
    fabric_llpp0_bvalid_s_i                      : in  std_logic;  -- dahlia_llpp0_bvalid_s_o
    fabric_llpp0_rdata_s_i1                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i2                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i3                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i4                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i5                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i6                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i7                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i8                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i9                      : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i10                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i11                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i12                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i13                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i14                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i15                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i16                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i17                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i18                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i19                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i20                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i21                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i22                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i23                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i24                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i25                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i26                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i27                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i28                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i29                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i30                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i31                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rdata_s_i32                     : in  std_logic;  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rid_s_i1                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i2                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i3                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i4                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i5                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i6                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i7                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i8                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i9                        : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i10                       : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i11                       : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rid_s_i12                       : in  std_logic;  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rlast_s_i                       : in  std_logic;  -- dahlia_llpp0_rlast_s_o
    fabric_llpp0_rresp_s_i1                      : in  std_logic;  -- dahlia_llpp0_rresp_s_o
    fabric_llpp0_rresp_s_i2                      : in  std_logic;  -- dahlia_llpp0_rresp_s_o
    fabric_llpp0_rvalid_s_i                      : in  std_logic;  -- dahlia_llpp0_rvalid_s_o
    fabric_llpp0_wready_s_i                      : in  std_logic;  -- dahlia_llpp0_wready_s_o
    fabric_llpp1_araddr_s_o1                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o2                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o3                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o4                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o5                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o6                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o7                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o8                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o9                     : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o10                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o11                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o12                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o13                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o14                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o15                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o16                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o17                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o18                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o19                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o20                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o21                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o22                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o23                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o24                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o25                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o26                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o27                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o28                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o29                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o30                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o31                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_araddr_s_o32                    : out std_logic;  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_arburst_s_o1                    : out std_logic;  -- dahlia_llpp1_arburst_s_i
    fabric_llpp1_arburst_s_o2                    : out std_logic;  -- dahlia_llpp1_arburst_s_i
    fabric_llpp1_arcache_s_o1                    : out std_logic;  -- dahlia_llpp1_arcache_s_i
    fabric_llpp1_arcache_s_o2                    : out std_logic;  -- dahlia_llpp1_arcache_s_i
    fabric_llpp1_arcache_s_o3                    : out std_logic;  -- dahlia_llpp1_arcache_s_i
    fabric_llpp1_arcache_s_o4                    : out std_logic;  -- dahlia_llpp1_arcache_s_i
    fabric_llpp1_arid_s_o1                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o2                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o3                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o4                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o5                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o6                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o7                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o8                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o9                       : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o10                      : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o11                      : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arid_s_o12                      : out std_logic;  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arlen_s_o1                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o2                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o3                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o4                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o5                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o6                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o7                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlen_s_o8                      : out std_logic;  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlock_s_o                      : out std_logic;  -- dahlia_llpp1_arlock_s_i
    fabric_llpp1_arprot_s_o1                     : out std_logic;  -- dahlia_llpp1_arprot_s_i
    fabric_llpp1_arprot_s_o2                     : out std_logic;  -- dahlia_llpp1_arprot_s_i
    fabric_llpp1_arprot_s_o3                     : out std_logic;  -- dahlia_llpp1_arprot_s_i
    fabric_llpp1_arqos_s1_o1                     : out std_logic;  -- dahlia_llpp1_arqos_s1_i
    fabric_llpp1_arqos_s1_o2                     : out std_logic;  -- dahlia_llpp1_arqos_s1_i
    fabric_llpp1_arqos_s1_o3                     : out std_logic;  -- dahlia_llpp1_arqos_s1_i
    fabric_llpp1_arqos_s1_o4                     : out std_logic;  -- dahlia_llpp1_arqos_s1_i
    fabric_llpp1_arsize_s_o1                     : out std_logic;  -- dahlia_llpp1_arsize_s_i
    fabric_llpp1_arsize_s_o2                     : out std_logic;  -- dahlia_llpp1_arsize_s_i
    fabric_llpp1_arsize_s_o3                     : out std_logic;  -- dahlia_llpp1_arsize_s_i
    fabric_llpp1_arvalid_s_o                     : out std_logic;  -- dahlia_llpp1_arvalid_s_i
    fabric_llpp1_awaddr_s_o1                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o2                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o3                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o4                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o5                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o6                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o7                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o8                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o9                     : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o10                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o11                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o12                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o13                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o14                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o15                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o16                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o17                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o18                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o19                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o20                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o21                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o22                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o23                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o24                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o25                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o26                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o27                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o28                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o29                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o30                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o31                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awaddr_s_o32                    : out std_logic;  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awburst_s_o1                    : out std_logic;  -- dahlia_llpp1_awburst_s_i
    fabric_llpp1_awburst_s_o2                    : out std_logic;  -- dahlia_llpp1_awburst_s_i
    fabric_llpp1_awcache_s_o1                    : out std_logic;  -- dahlia_llpp1_awcache_s_i
    fabric_llpp1_awcache_s_o2                    : out std_logic;  -- dahlia_llpp1_awcache_s_i
    fabric_llpp1_awcache_s_o3                    : out std_logic;  -- dahlia_llpp1_awcache_s_i
    fabric_llpp1_awcache_s_o4                    : out std_logic;  -- dahlia_llpp1_awcache_s_i
    fabric_llpp1_awid_s_o1                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o2                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o3                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o4                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o5                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o6                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o7                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o8                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o9                       : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o10                      : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o11                      : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awid_s_o12                      : out std_logic;  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awlen_s_o1                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o2                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o3                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o4                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o5                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o6                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o7                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlen_s_o8                      : out std_logic;  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlock_s_o                      : out std_logic;  -- dahlia_llpp1_awlock_s_i
    fabric_llpp1_awprot_s_o1                     : out std_logic;  -- dahlia_llpp1_awprot_s_i
    fabric_llpp1_awprot_s_o2                     : out std_logic;  -- dahlia_llpp1_awprot_s_i
    fabric_llpp1_awprot_s_o3                     : out std_logic;  -- dahlia_llpp1_awprot_s_i
    fabric_llpp1_awqos_s_o1                      : out std_logic;  -- dahlia_llpp1_awqos_s_i
    fabric_llpp1_awqos_s_o2                      : out std_logic;  -- dahlia_llpp1_awqos_s_i
    fabric_llpp1_awqos_s_o3                      : out std_logic;  -- dahlia_llpp1_awqos_s_i
    fabric_llpp1_awqos_s_o4                      : out std_logic;  -- dahlia_llpp1_awqos_s_i
    fabric_llpp1_awsize_s_o1                     : out std_logic;  -- dahlia_llpp1_awsize_s_i
    fabric_llpp1_awsize_s_o2                     : out std_logic;  -- dahlia_llpp1_awsize_s_i
    fabric_llpp1_awsize_s_o3                     : out std_logic;  -- dahlia_llpp1_awsize_s_i
    fabric_llpp1_awvalid_s_o                     : out std_logic;  -- dahlia_llpp1_awvalid_s_i
    fabric_llpp1_bready_s_o                      : out std_logic;  -- dahlia_llpp1_bready_s_i
    fabric_llpp1_rready_s_o                      : out std_logic;  -- dahlia_llpp1_rready_s_i
    fabric_llpp1_wdata_s_o1                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o2                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o3                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o4                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o5                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o6                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o7                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o8                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o9                      : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o10                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o11                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o12                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o13                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o14                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o15                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o16                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o17                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o18                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o19                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o20                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o21                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o22                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o23                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o24                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o25                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o26                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o27                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o28                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o29                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o30                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o31                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wdata_s_o32                     : out std_logic;  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wlast_s_o                       : out std_logic;  -- dahlia_llpp1_wlast_s_i
    fabric_llpp1_wstrb_s_o1                      : out std_logic;  -- dahlia_llpp1_wstrb_s_i
    fabric_llpp1_wstrb_s_o2                      : out std_logic;  -- dahlia_llpp1_wstrb_s_i
    fabric_llpp1_wstrb_s_o3                      : out std_logic;  -- dahlia_llpp1_wstrb_s_i
    fabric_llpp1_wstrb_s_o4                      : out std_logic;  -- dahlia_llpp1_wstrb_s_i
    fabric_llpp1_wvalid_s_o                      : out std_logic;  -- dahlia_llpp1_wvalid_s_i
    fabric_llpp1_arready_s_i                     : in  std_logic;  -- dahlia_llpp1_arready_s_o
    fabric_llpp1_awready_s_i                     : in  std_logic;  -- dahlia_llpp1_awready_s_o
    fabric_llpp1_bid_s_i1                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i2                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i3                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i4                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i5                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i6                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i7                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i8                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i9                        : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i10                       : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i11                       : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bid_s_i12                       : in  std_logic;  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bresp_s_i1                      : in  std_logic;  -- dahlia_llpp1_bresp_s_o
    fabric_llpp1_bresp_s_i2                      : in  std_logic;  -- dahlia_llpp1_bresp_s_o
    fabric_llpp1_bvalid_s_i                      : in  std_logic;  -- dahlia_llpp1_bvalid_s_o
    fabric_llpp1_rdata_s_i1                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i2                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i3                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i4                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i5                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i6                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i7                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i8                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i9                      : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i10                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i11                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i12                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i13                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i14                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i15                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i16                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i17                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i18                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i19                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i20                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i21                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i22                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i23                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i24                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i25                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i26                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i27                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i28                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i29                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i30                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i31                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rdata_s_i32                     : in  std_logic;  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rid_s_i1                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i2                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i3                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i4                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i5                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i6                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i7                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i8                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i9                        : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i10                       : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i11                       : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rid_s_i12                       : in  std_logic;  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rlast_s_i                       : in  std_logic;  -- dahlia_llpp1_rlast_s_o
    fabric_llpp1_rresp_s_i1                      : in  std_logic;  -- dahlia_llpp1_rresp_s_o
    fabric_llpp1_rresp_s_i2                      : in  std_logic;  -- dahlia_llpp1_rresp_s_o
    fabric_llpp1_rvalid_s_i                      : in  std_logic;  -- dahlia_llpp1_rvalid_s_o
    fabric_llpp1_wready_s_i                      : in  std_logic;  -- dahlia_llpp1_wready_s_o
    fabric_llpp2_araddr_s_o1                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o2                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o3                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o4                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o5                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o6                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o7                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o8                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o9                     : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o10                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o11                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o12                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o13                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o14                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o15                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o16                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o17                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o18                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o19                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o20                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o21                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o22                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o23                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o24                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o25                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o26                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o27                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o28                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o29                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o30                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o31                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_araddr_s_o32                    : out std_logic;  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_arburst_s_o1                    : out std_logic;  -- dahlia_llpp2_arburst_s_i
    fabric_llpp2_arburst_s_o2                    : out std_logic;  -- dahlia_llpp2_arburst_s_i
    fabric_llpp2_arcache_s_o1                    : out std_logic;  -- dahlia_llpp2_arcache_s_i
    fabric_llpp2_arcache_s_o2                    : out std_logic;  -- dahlia_llpp2_arcache_s_i
    fabric_llpp2_arcache_s_o3                    : out std_logic;  -- dahlia_llpp2_arcache_s_i
    fabric_llpp2_arcache_s_o4                    : out std_logic;  -- dahlia_llpp2_arcache_s_i
    fabric_llpp2_arid_s_o1                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o2                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o3                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o4                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o5                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o6                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o7                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o8                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o9                       : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o10                      : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o11                      : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arid_s_o12                      : out std_logic;  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arlen_s_o1                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o2                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o3                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o4                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o5                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o6                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o7                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlen_s_o8                      : out std_logic;  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlock_s_o                      : out std_logic;  -- dahlia_llpp2_arlock_s_i
    fabric_llpp2_arprot_s_o1                     : out std_logic;  -- dahlia_llpp2_arprot_s_i
    fabric_llpp2_arprot_s_o2                     : out std_logic;  -- dahlia_llpp2_arprot_s_i
    fabric_llpp2_arprot_s_o3                     : out std_logic;  -- dahlia_llpp2_arprot_s_i
    fabric_llpp2_arqos_s_o1                      : out std_logic;  -- dahlia_llpp2_arqos_s_i
    fabric_llpp2_arqos_s_o2                      : out std_logic;  -- dahlia_llpp2_arqos_s_i
    fabric_llpp2_arqos_s_o3                      : out std_logic;  -- dahlia_llpp2_arqos_s_i
    fabric_llpp2_arqos_s_o4                      : out std_logic;  -- dahlia_llpp2_arqos_s_i
    fabric_llpp2_arsize_s_o1                     : out std_logic;  -- dahlia_llpp2_arsize_s_i
    fabric_llpp2_arsize_s_o2                     : out std_logic;  -- dahlia_llpp2_arsize_s_i
    fabric_llpp2_arsize_s_o3                     : out std_logic;  -- dahlia_llpp2_arsize_s_i
    fabric_llpp2_arvalid_s_o                     : out std_logic;  -- dahlia_llpp2_arvalid_s_i
    fabric_llpp2_awaddr_s_o1                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o2                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o3                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o4                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o5                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o6                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o7                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o8                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o9                     : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o10                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o11                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o12                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o13                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o14                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o15                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o16                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o17                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o18                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o19                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o20                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o21                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o22                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o23                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o24                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o25                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o26                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o27                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o28                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o29                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o30                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o31                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awaddr_s_o32                    : out std_logic;  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awburst_s_o1                    : out std_logic;  -- dahlia_llpp2_awburst_s_i
    fabric_llpp2_awburst_s_o2                    : out std_logic;  -- dahlia_llpp2_awburst_s_i
    fabric_llpp2_awcache_s_o1                    : out std_logic;  -- dahlia_llpp2_awcache_s_i
    fabric_llpp2_awcache_s_o2                    : out std_logic;  -- dahlia_llpp2_awcache_s_i
    fabric_llpp2_awcache_s_o3                    : out std_logic;  -- dahlia_llpp2_awcache_s_i
    fabric_llpp2_awcache_s_o4                    : out std_logic;  -- dahlia_llpp2_awcache_s_i
    fabric_llpp2_awid_s_o1                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o2                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o3                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o4                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o5                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o6                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o7                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o8                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o9                       : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o10                      : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o11                      : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awid_s_o12                      : out std_logic;  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awlen_s_o1                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o2                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o3                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o4                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o5                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o6                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o7                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlen_s_o8                      : out std_logic;  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlock_s_o                      : out std_logic;  -- dahlia_llpp2_awlock_s_i
    fabric_llpp2_awprot_s_o1                     : out std_logic;  -- dahlia_llpp2_awprot_s_i
    fabric_llpp2_awprot_s_o2                     : out std_logic;  -- dahlia_llpp2_awprot_s_i
    fabric_llpp2_awprot_s_o3                     : out std_logic;  -- dahlia_llpp2_awprot_s_i
    fabric_llpp2_awqos_s_o1                      : out std_logic;  -- dahlia_llpp2_awqos_s_i
    fabric_llpp2_awqos_s_o2                      : out std_logic;  -- dahlia_llpp2_awqos_s_i
    fabric_llpp2_awqos_s_o3                      : out std_logic;  -- dahlia_llpp2_awqos_s_i
    fabric_llpp2_awqos_s_o4                      : out std_logic;  -- dahlia_llpp2_awqos_s_i
    fabric_llpp2_awsize_s_o1                     : out std_logic;  -- dahlia_llpp2_awsize_s_i
    fabric_llpp2_awsize_s_o2                     : out std_logic;  -- dahlia_llpp2_awsize_s_i
    fabric_llpp2_awsize_s_o3                     : out std_logic;  -- dahlia_llpp2_awsize_s_i
    fabric_llpp2_awvalid_s_o                     : out std_logic;  -- dahlia_llpp2_awvalid_s_i
    fabric_llpp2_bready_s_o                      : out std_logic;  -- dahlia_llpp2_bready_s_i
    fabric_llpp2_rready_s_o                      : out std_logic;  -- dahlia_llpp2_rready_s_i
    fabric_llpp2_wdata_s_o1                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o2                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o3                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o4                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o5                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o6                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o7                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o8                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o9                      : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o10                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o11                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o12                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o13                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o14                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o15                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o16                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o17                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o18                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o19                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o20                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o21                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o22                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o23                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o24                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o25                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o26                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o27                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o28                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o29                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o30                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o31                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wdata_s_o32                     : out std_logic;  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wlast_s_o                       : out std_logic;  -- dahlia_llpp2_wlast_s_i
    fabric_llpp2_wstrb_s_o1                      : out std_logic;  -- dahlia_llpp2_wstrb_s_i
    fabric_llpp2_wstrb_s_o2                      : out std_logic;  -- dahlia_llpp2_wstrb_s_i
    fabric_llpp2_wstrb_s_o3                      : out std_logic;  -- dahlia_llpp2_wstrb_s_i
    fabric_llpp2_wstrb_s_o4                      : out std_logic;  -- dahlia_llpp2_wstrb_s_i
    fabric_llpp2_wvalid_s_o                      : out std_logic;  -- dahlia_llpp2_wvalid_s_i
    fabric_llpp2_arready_s_i                     : in  std_logic;  -- dahlia_llpp2_arready_s_o
    fabric_llpp2_awready_s_i                     : in  std_logic;  -- dahlia_llpp2_awready_s_o
    fabric_llpp2_bid_s_i1                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i2                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i3                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i4                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i5                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i6                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i7                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i8                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i9                        : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i10                       : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i11                       : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bid_s_i12                       : in  std_logic;  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bresp_s_i1                      : in  std_logic;  -- dahlia_llpp2_bresp_s_o
    fabric_llpp2_bresp_s_i2                      : in  std_logic;  -- dahlia_llpp2_bresp_s_o
    fabric_llpp2_bvalid_s_i                      : in  std_logic;  -- dahlia_llpp2_bvalid_s_o
    fabric_llpp2_rdata_s_i1                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i2                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i3                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i4                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i5                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i6                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i7                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i8                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i9                      : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i10                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i11                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i12                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i13                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i14                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i15                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i16                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i17                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i18                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i19                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i20                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i21                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i22                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i23                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i24                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i25                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i26                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i27                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i28                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i29                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i30                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i31                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rdata_s_i32                     : in  std_logic;  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rid_s_i1                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i2                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i3                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i4                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i5                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i6                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i7                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i8                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i9                        : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i10                       : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i11                       : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rid_s_i12                       : in  std_logic;  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rlast_s_i                       : in  std_logic;  -- dahlia_llpp2_rlast_s_o
    fabric_llpp2_rresp_s_i1                      : in  std_logic;  -- dahlia_llpp2_rresp_s_o
    fabric_llpp2_rresp_s_i2                      : in  std_logic;  -- dahlia_llpp2_rresp_s_o
    fabric_llpp2_rvalid_s_i                      : in  std_logic;  -- dahlia_llpp2_rvalid_s_o
    fabric_llpp2_wready_s_i                      : in  std_logic;  -- dahlia_llpp2_wready_s_o
    fabric_llpp3_araddr_s_o1                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o2                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o3                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o4                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o5                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o6                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o7                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o8                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o9                     : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o10                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o11                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o12                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o13                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o14                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o15                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o16                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o17                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o18                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o19                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o20                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o21                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o22                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o23                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o24                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o25                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o26                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o27                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o28                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o29                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o30                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o31                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_araddr_s_o32                    : out std_logic;  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_arburst_s_o1                    : out std_logic;  -- dahlia_llpp3_arburst_s_i
    fabric_llpp3_arburst_s_o2                    : out std_logic;  -- dahlia_llpp3_arburst_s_i
    fabric_llpp3_arcache_s_o1                    : out std_logic;  -- dahlia_llpp3_arcache_s_i
    fabric_llpp3_arcache_s_o2                    : out std_logic;  -- dahlia_llpp3_arcache_s_i
    fabric_llpp3_arcache_s_o3                    : out std_logic;  -- dahlia_llpp3_arcache_s_i
    fabric_llpp3_arcache_s_o4                    : out std_logic;  -- dahlia_llpp3_arcache_s_i
    fabric_llpp3_arid_s_o1                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o2                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o3                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o4                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o5                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o6                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o7                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o8                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o9                       : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o10                      : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o11                      : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arid_s_o12                      : out std_logic;  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arlen_s_o1                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o2                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o3                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o4                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o5                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o6                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o7                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlen_s_o8                      : out std_logic;  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlock_s_o                      : out std_logic;  -- dahlia_llpp3_arlock_s_i
    fabric_llpp3_arprot_s_o1                     : out std_logic;  -- dahlia_llpp3_arprot_s_i
    fabric_llpp3_arprot_s_o2                     : out std_logic;  -- dahlia_llpp3_arprot_s_i
    fabric_llpp3_arprot_s_o3                     : out std_logic;  -- dahlia_llpp3_arprot_s_i
    fabric_llpp3_arqos_s_o1                      : out std_logic;  -- dahlia_llpp3_arqos_s_i
    fabric_llpp3_arqos_s_o2                      : out std_logic;  -- dahlia_llpp3_arqos_s_i
    fabric_llpp3_arqos_s_o3                      : out std_logic;  -- dahlia_llpp3_arqos_s_i
    fabric_llpp3_arqos_s_o4                      : out std_logic;  -- dahlia_llpp3_arqos_s_i
    fabric_llpp3_arsize_s_o1                     : out std_logic;  -- dahlia_llpp3_arsize_s_i
    fabric_llpp3_arsize_s_o2                     : out std_logic;  -- dahlia_llpp3_arsize_s_i
    fabric_llpp3_arsize_s_o3                     : out std_logic;  -- dahlia_llpp3_arsize_s_i
    fabric_llpp3_arvalid_s_o                     : out std_logic;  -- dahlia_llpp3_arvalid_s_i
    fabric_llpp3_awaddr_s_o1                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o2                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o3                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o4                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o5                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o6                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o7                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o8                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o9                     : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o10                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o11                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o12                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o13                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o14                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o15                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o16                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o17                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o18                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o19                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o20                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o21                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o22                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o23                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o24                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o25                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o26                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o27                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o28                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o29                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o30                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o31                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awaddr_s_o32                    : out std_logic;  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awburst_s_o1                    : out std_logic;  -- dahlia_llpp3_awburst_s_i
    fabric_llpp3_awburst_s_o2                    : out std_logic;  -- dahlia_llpp3_awburst_s_i
    fabric_llpp3_awcache_s_o1                    : out std_logic;  -- dahlia_llpp3_awcache_s_i
    fabric_llpp3_awcache_s_o2                    : out std_logic;  -- dahlia_llpp3_awcache_s_i
    fabric_llpp3_awcache_s_o3                    : out std_logic;  -- dahlia_llpp3_awcache_s_i
    fabric_llpp3_awcache_s_o4                    : out std_logic;  -- dahlia_llpp3_awcache_s_i
    fabric_llpp3_awid_s_o1                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o2                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o3                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o4                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o5                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o6                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o7                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o8                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o9                       : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o10                      : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o11                      : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awid_s_o12                      : out std_logic;  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awlen_s_o1                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o2                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o3                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o4                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o5                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o6                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o7                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlen_s_o8                      : out std_logic;  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlock_s_o                      : out std_logic;  -- dahlia_llpp3_awlock_s_i
    fabric_llpp3_awprot_s_o1                     : out std_logic;  -- dahlia_llpp3_awprot_s_i
    fabric_llpp3_awprot_s_o2                     : out std_logic;  -- dahlia_llpp3_awprot_s_i
    fabric_llpp3_awprot_s_o3                     : out std_logic;  -- dahlia_llpp3_awprot_s_i
    fabric_llpp3_awqos_s_o1                      : out std_logic;  -- dahlia_llpp3_awqos_s_i
    fabric_llpp3_awqos_s_o2                      : out std_logic;  -- dahlia_llpp3_awqos_s_i
    fabric_llpp3_awqos_s_o3                      : out std_logic;  -- dahlia_llpp3_awqos_s_i
    fabric_llpp3_awqos_s_o4                      : out std_logic;  -- dahlia_llpp3_awqos_s_i
    fabric_llpp3_awsize_s_o1                     : out std_logic;  -- dahlia_llpp3_awsize_s_i
    fabric_llpp3_awsize_s_o2                     : out std_logic;  -- dahlia_llpp3_awsize_s_i
    fabric_llpp3_awsize_s_o3                     : out std_logic;  -- dahlia_llpp3_awsize_s_i
    fabric_llpp3_awvalid_s_o                     : out std_logic;  -- dahlia_llpp3_awvalid_s_i
    fabric_llpp3_bready_s_o                      : out std_logic;  -- dahlia_llpp3_bready_s_i
    fabric_llpp3_rready_s_o                      : out std_logic;  -- dahlia_llpp3_rready_s_i
    fabric_llpp3_wdata_s_o1                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o2                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o3                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o4                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o5                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o6                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o7                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o8                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o9                      : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o10                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o11                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o12                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o13                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o14                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o15                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o16                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o17                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o18                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o19                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o20                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o21                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o22                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o23                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o24                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o25                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o26                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o27                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o28                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o29                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o30                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o31                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wdata_s_o32                     : out std_logic;  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wlast_s_o                       : out std_logic;  -- dahlia_llpp3_wlast_s_i
    fabric_llpp3_wstrb_s_o1                      : out std_logic;  -- dahlia_llpp3_wstrb_s_i
    fabric_llpp3_wstrb_s_o2                      : out std_logic;  -- dahlia_llpp3_wstrb_s_i
    fabric_llpp3_wstrb_s_o3                      : out std_logic;  -- dahlia_llpp3_wstrb_s_i
    fabric_llpp3_wstrb_s_o4                      : out std_logic;  -- dahlia_llpp3_wstrb_s_i
    fabric_llpp3_wvalid_s_o                      : out std_logic;  -- dahlia_llpp3_wvalid_s_i
    fabric_llpp3_arready_s_i                     : in  std_logic;  -- dahlia_llpp3_arready_s_o
    fabric_llpp3_awready_s_i                     : in  std_logic;  -- dahlia_llpp3_awready_s_o
    fabric_llpp3_bid_s_i1                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i2                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i3                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i4                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i5                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i6                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i7                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i8                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i9                        : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i10                       : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i11                       : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bid_s_i12                       : in  std_logic;  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bresp_s_i1                      : in  std_logic;  -- dahlia_llpp3_bresp_s_o
    fabric_llpp3_bresp_s_i2                      : in  std_logic;  -- dahlia_llpp3_bresp_s_o
    fabric_llpp3_bvalid_s_i                      : in  std_logic;  -- dahlia_llpp3_bvalid_s_o
    fabric_llpp3_rdata_s_i1                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i2                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i3                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i4                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i5                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i6                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i7                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i8                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i9                      : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i10                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i11                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i12                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i13                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i14                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i15                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i16                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i17                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i18                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i19                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i20                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i21                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i22                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i23                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i24                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i25                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i26                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i27                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i28                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i29                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i30                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i31                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rdata_s_i32                     : in  std_logic;  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rid_s_i1                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i2                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i3                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i4                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i5                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i6                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i7                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i8                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i9                        : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i10                       : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i11                       : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rid_s_i12                       : in  std_logic;  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rlast_s_i                       : in  std_logic;  -- dahlia_llpp3_rlast_s_o
    fabric_llpp3_rresp_s_i1                      : in  std_logic;  -- dahlia_llpp3_rresp_s_o
    fabric_llpp3_rresp_s_i2                      : in  std_logic;  -- dahlia_llpp3_rresp_s_o
    fabric_llpp3_rvalid_s_i                      : in  std_logic;  -- dahlia_llpp3_rvalid_s_o
    fabric_llpp3_wready_s_i                      : in  std_logic;  -- dahlia_llpp3_wready_s_o
    fabric_qos_pprdata_o1                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o2                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o3                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o4                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o5                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o6                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o7                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o8                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o9                        : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o10                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o11                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o12                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o13                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o14                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o15                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o16                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o17                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o18                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o19                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o20                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o21                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o22                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o23                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o24                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o25                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o26                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o27                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o28                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o29                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o30                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o31                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_pprdata_o32                       : out std_logic;  -- dahlia_qos_pprdata_i
    fabric_qos_ppready_o                         : out std_logic;  -- dahlia_qos_ppready_i
    fabric_qos_ppslverr_o                        : out std_logic;  -- dahlia_qos_ppslverr_i
    fabric_qos_pclk_i                            : in  std_logic;  -- dahlia_qos_pclk_o
    fabric_qos_ppaddr_i1                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i2                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i3                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i4                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i5                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i6                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i7                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i8                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i9                         : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i10                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i11                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i12                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i13                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i14                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i15                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i16                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i17                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i18                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i19                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i20                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i21                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i22                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i23                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i24                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i25                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i26                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i27                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i28                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i29                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i30                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i31                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppaddr_i32                        : in  std_logic;  -- dahlia_qos_ppaddr_o
    fabric_qos_ppenable_i                        : in  std_logic;  -- dahlia_qos_ppenable_o
    fabric_qos_ppwdata_i1                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i2                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i3                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i4                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i5                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i6                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i7                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i8                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i9                        : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i10                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i11                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i12                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i13                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i14                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i15                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i16                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i17                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i18                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i19                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i20                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i21                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i22                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i23                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i24                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i25                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i26                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i27                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i28                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i29                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i30                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i31                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwdata_i32                       : in  std_logic;  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwrite_i                         : in  std_logic;  -- dahlia_qos_ppwrite_o
    fabric_qos_presetn_i                         : in  std_logic;  -- dahlia_qos_presetn_o
    fabric_qos_psel_i                            : in  std_logic;  -- dahlia_qos_psel_o
    fabric_tnd_hssl_flushin_o                    : out std_logic;  -- dahlia_tnd_hssl_flushin_i
    fabric_tnd_hssl_trigin_o                     : out std_logic;  -- dahlia_tnd_hssl_trigin_i
    fabric_tnd_fpga_apb_master_paddr_o1          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o2          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o3          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o4          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o5          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o6          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o7          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o8          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o9          : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o10         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o11         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o12         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o13         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o14         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o15         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o16         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o17         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o18         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o19         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o20         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o21         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o22         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o23         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o24         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o25         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o26         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o27         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o28         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o29         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o30         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o31         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_paddr_o32         : out std_logic;  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_penable_o         : out std_logic;  -- dahlia_tnd_fpga_apb_master_penable_i
    fabric_tnd_fpga_apb_master_psel_o            : out std_logic;  -- dahlia_tnd_fpga_apb_master_psel_i
    fabric_tnd_fpga_apb_master_pwdata_o1         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o2         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o3         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o4         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o5         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o6         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o7         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o8         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o9         : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o10        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o11        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o12        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o13        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o14        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o15        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o16        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o17        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o18        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o19        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o20        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o21        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o22        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o23        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o24        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o25        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o26        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o27        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o28        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o29        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o30        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o31        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwdata_o32        : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwrite_o          : out std_logic;  -- dahlia_tnd_fpga_apb_master_pwrite_i
    fabric_tnd_fpga_atb_master_afvalid_o         : out std_logic;  -- dahlia_tnd_fpga_atb_master_afvalid_i
    fabric_tnd_fpga_atb_master_atready_o         : out std_logic;  -- dahlia_tnd_fpga_atb_master_atready_i
    fabric_tnd_fpga_atb_master_syncreq_o         : out std_logic;  -- dahlia_tnd_fpga_atb_master_syncreq_i
    fabric_tnd_hssl_apb_master_paddr_o1          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o2          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o3          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o4          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o5          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o6          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o7          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o8          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o9          : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o10         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o11         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o12         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o13         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o14         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o15         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o16         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o17         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o18         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o19         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o20         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o21         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o22         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o23         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o24         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o25         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o26         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o27         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o28         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o29         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o30         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o31         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_paddr_o32         : out std_logic;  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_penable_o         : out std_logic;  -- dahlia_tnd_hssl_apb_master_penable_i
    fabric_tnd_hssl_apb_master_psel_o            : out std_logic;  -- dahlia_tnd_hssl_apb_master_psel_i
    fabric_tnd_hssl_apb_master_pwdata_o1         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o2         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o3         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o4         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o5         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o6         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o7         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o8         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o9         : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o10        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o11        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o12        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o13        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o14        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o15        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o16        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o17        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o18        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o19        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o20        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o21        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o22        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o23        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o24        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o25        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o26        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o27        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o28        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o29        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o30        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o31        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwdata_o32        : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwrite_o          : out std_logic;  -- dahlia_tnd_hssl_apb_master_pwrite_i
    fabric_tnd_hssl_atb_master_afready_o         : out std_logic;  -- dahlia_tnd_hssl_atb_master_afready_i
    fabric_tnd_hssl_atb_master_atbytes_o1        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atbytes_i
    fabric_tnd_hssl_atb_master_atbytes_o2        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atbytes_i
    fabric_tnd_hssl_atb_master_atbytes_o3        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atbytes_i
    fabric_tnd_hssl_atb_master_atbytes_o4        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atbytes_i
    fabric_tnd_hssl_atb_master_atdata_o1         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o2         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o3         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o4         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o5         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o6         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o7         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o8         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o9         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o10        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o11        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o12        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o13        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o14        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o15        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o16        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o17        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o18        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o19        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o20        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o21        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o22        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o23        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o24        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o25        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o26        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o27        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o28        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o29        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o30        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o31        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o32        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o33        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o34        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o35        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o36        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o37        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o38        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o39        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o40        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o41        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o42        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o43        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o44        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o45        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o46        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o47        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o48        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o49        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o50        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o51        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o52        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o53        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o54        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o55        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o56        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o57        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o58        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o59        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o60        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o61        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o62        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o63        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o64        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o65        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o66        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o67        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o68        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o69        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o70        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o71        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o72        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o73        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o74        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o75        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o76        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o77        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o78        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o79        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o80        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o81        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o82        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o83        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o84        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o85        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o86        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o87        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o88        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o89        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o90        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o91        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o92        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o93        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o94        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o95        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o96        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o97        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o98        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o99        : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o100       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o101       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o102       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o103       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o104       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o105       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o106       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o107       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o108       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o109       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o110       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o111       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o112       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o113       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o114       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o115       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o116       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o117       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o118       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o119       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o120       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o121       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o122       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o123       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o124       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o125       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o126       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o127       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atdata_o128       : out std_logic;  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atid_o1           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o2           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o3           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o4           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o5           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o6           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atid_o7           : out std_logic;  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atvalid_o         : out std_logic;  -- dahlia_tnd_hssl_atb_master_atvalid_i
    fabric_tnd_trace_clk_traceoutportintf_o      : out std_logic;  -- dahlia_tnd_trace_clk_traceoutportintf_i
    fabric_tnd_trace_ctl_traceoutportintf_o      : out std_logic;  -- dahlia_tnd_trace_ctl_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o1    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o2    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o3    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o4    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o5    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o6    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o7    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o8    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o9    : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o10   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o11   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o12   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o13   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o14   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o15   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o16   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o17   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o18   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o19   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o20   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o21   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o22   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o23   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o24   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o25   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o26   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o27   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o28   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o29   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o30   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o31   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o32   : out std_logic;  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tsvalue_tsgen_fpga_o1                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o2                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o3                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o4                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o5                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o6                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o7                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o8                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o9                 : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o10                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o11                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o12                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o13                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o14                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o15                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o16                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o17                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o18                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o19                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o20                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o21                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o22                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o23                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o24                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o25                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o26                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o27                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o28                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o29                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o30                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o31                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o32                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o33                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o34                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o35                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o36                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o37                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o38                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o39                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o40                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o41                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o42                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o43                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o44                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o45                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o46                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o47                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o48                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o49                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o50                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o51                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o52                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o53                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o54                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o55                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o56                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o57                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o58                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o59                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o60                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o61                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o62                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o63                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tsvalue_tsgen_fpga_o64                : out std_logic;  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tnd_fpga_apb_master_prdata_i1         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i2         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i3         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i4         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i5         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i6         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i7         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i8         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i9         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i10        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i11        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i12        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i13        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i14        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i15        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i16        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i17        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i18        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i19        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i20        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i21        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i22        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i23        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i24        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i25        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i26        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i27        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i28        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i29        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i30        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i31        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_prdata_i32        : in  std_logic;  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_pready_i          : in  std_logic;  -- dahlia_tnd_fpga_apb_master_pready_o
    fabric_tnd_fpga_apb_master_pslverr_i         : in  std_logic;  -- dahlia_tnd_fpga_apb_master_pslverr_o
    fabric_tnd_fpga_atb_master_afready_i         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_afready_o
    fabric_tnd_fpga_atb_master_atbytes_i1        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atbytes_o
    fabric_tnd_fpga_atb_master_atbytes_i2        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atbytes_o
    fabric_tnd_fpga_atb_master_atbytes_i3        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atbytes_o
    fabric_tnd_fpga_atb_master_atbytes_i4        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atbytes_o
    fabric_tnd_fpga_atb_master_atdata_i1         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i2         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i3         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i4         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i5         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i6         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i7         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i8         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i9         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i10        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i11        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i12        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i13        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i14        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i15        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i16        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i17        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i18        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i19        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i20        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i21        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i22        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i23        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i24        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i25        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i26        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i27        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i28        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i29        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i30        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i31        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i32        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i33        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i34        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i35        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i36        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i37        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i38        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i39        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i40        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i41        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i42        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i43        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i44        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i45        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i46        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i47        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i48        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i49        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i50        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i51        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i52        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i53        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i54        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i55        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i56        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i57        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i58        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i59        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i60        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i61        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i62        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i63        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i64        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i65        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i66        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i67        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i68        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i69        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i70        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i71        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i72        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i73        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i74        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i75        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i76        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i77        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i78        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i79        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i80        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i81        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i82        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i83        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i84        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i85        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i86        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i87        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i88        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i89        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i90        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i91        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i92        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i93        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i94        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i95        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i96        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i97        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i98        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i99        : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i100       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i101       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i102       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i103       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i104       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i105       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i106       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i107       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i108       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i109       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i110       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i111       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i112       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i113       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i114       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i115       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i116       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i117       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i118       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i119       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i120       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i121       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i122       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i123       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i124       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i125       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i126       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i127       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atdata_i128       : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atid_i1           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i2           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i3           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i4           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i5           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i6           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atid_i7           : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atvalid_i         : in  std_logic;  -- dahlia_tnd_fpga_atb_master_atvalid_o
    fabric_tnd_hssl_apb_master_prdata_i1         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i2         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i3         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i4         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i5         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i6         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i7         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i8         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i9         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i10        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i11        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i12        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i13        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i14        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i15        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i16        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i17        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i18        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i19        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i20        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i21        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i22        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i23        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i24        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i25        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i26        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i27        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i28        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i29        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i30        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i31        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_prdata_i32        : in  std_logic;  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_pready_i          : in  std_logic;  -- dahlia_tnd_hssl_apb_master_pready_o
    fabric_tnd_hssl_apb_master_pslverr_i         : in  std_logic;  -- dahlia_tnd_hssl_apb_master_pslverr_o
    fabric_tnd_hssl_atb_master_afvalid_i         : in  std_logic;  -- dahlia_tnd_hssl_atb_master_afvalid_o
    fabric_tnd_hssl_atb_master_atready_i         : in  std_logic;  -- dahlia_tnd_hssl_atb_master_atready_o
    fabric_tnd_hssl_atb_master_syncreq_i         : in  std_logic;  -- dahlia_tnd_hssl_atb_master_syncreq_o
    fabric_watchdog0_signal_0_o                    : out std_logic;  -- dahlia_watchdog0_signal_0_i
    fabric_watchdog0_signal_1_o                    : out std_logic;  -- dahlia_watchdog0_signal_1_i
    fabric_watchdog1_signal_0_o                    : out std_logic;  -- dahlia_watchdog1_signal_0_i
    fabric_watchdog1_signal_1_o                    : out std_logic;  -- dahlia_watchdog1_signal_1_i
    fabric_watchdog2_signal_0_o                    : out std_logic;  -- dahlia_watchdog2_signal_0_i
    fabric_watchdog2_signal_1_o                    : out std_logic;  -- dahlia_watchdog2_signal_1_i
    fabric_watchdog3_signal_0_o                    : out std_logic;  -- dahlia_watchdog3_signal_0_i
    fabric_watchdog3_signal_1_o                    : out std_logic;  -- dahlia_watchdog3_signal_1_i
    fabric_tst_pll_lock_o1                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o2                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o3                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o4                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o5                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o6                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_tst_pll_lock_o7                       : out std_logic;  -- dahlia_tst_pll_lock_i
    fabric_soc_mon_sensor_alarm_o                : out std_logic;  -- dahlia_soc_mon_sensor_alarm_i
    fabric_erom_fpga_cpu0_dbgen_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu0_dbgen_o
    fabric_erom_fpga_cpu0_hiden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu0_hiden_o
    fabric_erom_fpga_cpu0_hniden_i               : in  std_logic;  -- dahlia_erom_fpga_cpu0_hniden_o
    fabric_erom_fpga_cpu0_niden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu0_niden_o
    fabric_erom_fpga_cpu1_dbgen_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu1_dbgen_o
    fabric_erom_fpga_cpu1_hiden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu1_hiden_o
    fabric_erom_fpga_cpu1_hniden_i               : in  std_logic;  -- dahlia_erom_fpga_cpu1_hniden_o
    fabric_erom_fpga_cpu1_niden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu1_niden_o
    fabric_erom_fpga_cpu2_dbgen_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu2_dbgen_o
    fabric_erom_fpga_cpu2_hiden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu2_hiden_o
    fabric_erom_fpga_cpu2_hniden_i               : in  std_logic;  -- dahlia_erom_fpga_cpu2_hniden_o
    fabric_erom_fpga_cpu2_niden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu2_niden_o
    fabric_erom_fpga_cpu3_dbgen_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu3_dbgen_o
    fabric_erom_fpga_cpu3_hiden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu3_hiden_o
    fabric_erom_fpga_cpu3_hniden_i               : in  std_logic;  -- dahlia_erom_fpga_cpu3_hniden_o
    fabric_erom_fpga_cpu3_niden_i                    : in  std_logic;  -- dahlia_erom_fpga_cpu3_niden_o
    fabric_erom_fpga_cs_dbgen_i                    : in  std_logic;  -- dahlia_erom_fpga_cs_dbgen_o
    fabric_erom_fpga_cs_niden_i                    : in  std_logic;  -- dahlia_erom_fpga_cs_niden_o
    fabric_erom_fpga_cs_deviceen_i               : in  std_logic;  -- dahlia_erom_fpga_cs_deviceen_o
    fabric_erom_fpga_cs_rst_n_i                    : in  std_logic;  -- dahlia_erom_fpga_cs_rst_n_o
    fabric_erom_fpga_debug_en_i                    : in  std_logic;  -- dahlia_erom_fpga_debug_en_o
    fabric_enable_TMR_i1                           : in  std_logic := '1';
    fabric_enable_TMR_i2                           : in  std_logic := '1';
    fabric_enable_TMR_i3                           : in  std_logic := '1'
);
end NX_SOC_INTERFACE;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--  NX_SOC_INTERFACE_WRAP definition
-- =================================================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library NX;
use NX.nxPackage.all;

entity NX_SOC_INTERFACE_WRAP is
generic (
    bsm_config : bit_vector(31 downto 0) := (others => '0');
    ahb_config : bit_vector(31 downto 0) := (others => '0')
);
port (
    -- dahlia <-> fabric
    fabric_lowskew_o                             : out std_logic_vector(1   downto 0);  -- dahlia_rstn_fpga_out_i / dahlia_clk_fpga_i
    fabric_lowskew_i                             : in  std_logic_vector(9   downto 0);  -- dahlia_clk_fpga_nic_o
    fabric_fpga_nic_rstn_i                       : in  std_logic_vector(9   downto 0);  -- dahlia_fpga_nic_rstn_o
    fabric_fpga_pmrstn_i                         : in  std_logic;                       -- dahlia_fpga_pmrstn_o
    fabric_fpga_sysrstn_i                        : in  std_logic;                       -- dahlia_fpga_sysrstn_o
    fabric_fpga_trigger_in_o                     : out std_logic_vector(7   downto 0);  -- dahlia_fpga_trigger_in_i
    fabric_fpga_trigger_out_i                    : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_trigger_out_o
    fabric_fpga_interrupt_in_i                   : in  std_logic_vector(119 downto 0);  -- dahlia_fpga_interrupt_in_o
    fabric_sysc_hold_on_debug_i                  : in  std_logic;                       -- dahlia_sysc_hold_on_debug_o
    fabric_fpga_events60_i                       : in  std_logic_vector(59  downto 0);  -- dahlia_fpga_events60_o
    fabric_fpga_araddr_axi_s1_o                  : out std_logic_vector(39  downto 0);  -- dahlia_fpga_araddr_axi_s1_i
    fabric_fpga_arburst_axi_s1_o                 : out std_logic_vector(1   downto 0);  -- dahlia_fpga_arburst_axi_s1_i
    fabric_fpga_arcache_axi_s1_o                 : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arcache_axi_s1_i
    fabric_fpga_arid_axi_s1_o                    : out std_logic_vector(11  downto 0);  -- dahlia_fpga_arid_axi_s1_i
    fabric_fpga_arlen_axi_s1_o                   : out std_logic_vector(7   downto 0);  -- dahlia_fpga_arlen_axi_s1_i
    fabric_fpga_arlock_axi_s1_o                  : out std_logic;                       -- dahlia_fpga_arlock_axi_s1_i
    fabric_fpga_arprot_axi_s1_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_arprot_axi_s1_i
    fabric_fpga_arqos_axi_s1_o                   : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arqos_axi_s1_i
    fabric_fpga_arregion_axi_s1_o                : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arregion_axi_s1_i
    fabric_fpga_arsize_axi_s1_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_arsize_axi_s1_i
    fabric_fpga_arvalid_axi_s1_o                 : out std_logic;                       -- dahlia_fpga_arvalid_axi_s1_i
    fabric_fpga_awaddr_axi_s1_o                  : out std_logic_vector(39  downto 0);  -- dahlia_fpga_awaddr_axi_s1_i
    fabric_fpga_awburst_axi_s1_o                 : out std_logic_vector(1   downto 0);  -- dahlia_fpga_awburst_axi_s1_i
    fabric_fpga_awcache_axi_s1_o                 : out std_logic_vector(3  downto 0);   -- dahlia_fpga_awcache_axi_s1_i
    fabric_fpga_awid_axi_s1_o                    : out std_logic_vector(11  downto 0);  -- dahlia_fpga_awid_axi_s1_i
    fabric_fpga_awlen_axi_s1_o                   : out std_logic_vector(7   downto 0);  -- dahlia_fpga_awlen_axi_s1_i
    fabric_fpga_awlock_axi_s1_o                  : out std_logic;                       -- dahlia_fpga_awlock_axi_s1_i
    fabric_fpga_awprot_axi_s1_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_awprot_axi_s1_i
    fabric_fpga_awqos_axi_s1_o                   : out std_logic_vector(3   downto 0);  -- dahlia_fpga_awqos_axi_s1_i
    fabric_fpga_awregion_axi_s1_o                : out std_logic_vector(3   downto 0);  -- dahlia_fpga_awregion_axi_s1_i
    fabric_fpga_awsize_axi_s1_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_awsize_axi_s1_i
    fabric_fpga_bready_axi_s1_o                  : out std_logic;                       -- dahlia_fpga_bready_axi_s1_i
    fabric_fpga_rready_axi_s1_o                  : out std_logic;                       -- dahlia_fpga_rready_axi_s1_i
    fabric_fpga_wdata_axi_s1_o                   : out std_logic_vector(127 downto 0);  -- dahlia_fpga_wdata_axi_s1_i
    fabric_fpga_wlast_axi_s1_o                   : out std_logic;                       -- dahlia_fpga_wlast_axi_s1_i
    fabric_fpga_wstrb_axi_s1_o                   : out std_logic_vector(15  downto 0);  -- dahlia_fpga_wstrb_axi_s1_i
    fabric_fpga_wvalid_axi_s1_o                  : out std_logic;                       -- dahlia_fpga_wvalid_axi_s1_i
    fabric_fpga_awvalid_axi_s1_o                 : out std_logic;                       -- dahlia_fpga_awvalid_axi_s1_i
    fabric_fpga_arready_axi_s1_i                 : in  std_logic;                       -- dahlia_fpga_arready_axi_s1_o
    fabric_fpga_awready_axi_s1_i                 : in  std_logic;                       -- dahlia_fpga_awready_axi_s1_o
    fabric_fpga_bid_axi_s1_i                     : in  std_logic_vector(11  downto 0);  -- dahlia_fpga_bid_axi_s1_o
    fabric_fpga_bresp_axi_s1_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_bresp_axi_s1_o
    fabric_fpga_bvalid_axi_s1_i                  : in  std_logic;                       -- dahlia_fpga_bvalid_axi_s1_o
    fabric_fpga_rdata_axi_s1_i                   : in  std_logic_vector(127 downto 0);  -- dahlia_fpga_rdata_axi_s1_o
    fabric_fpga_rid_axi_s1_i                     : in  std_logic_vector(11  downto 0);  -- dahlia_fpga_rid_axi_s1_o
    fabric_fpga_rlast_axi_s1_i                   : in  std_logic;                       -- dahlia_fpga_rlast_axi_s1_o
    fabric_fpga_rresp_axi_s1_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_rresp_axi_s1_o
    fabric_fpga_rvalid_axi_s1_i                  : in  std_logic;                       -- dahlia_fpga_rvalid_axi_s1_o
    fabric_fpga_wready_axi_s1_i                  : in  std_logic;                       -- dahlia_fpga_wready_axi_s1_o
    fabric_fpga_araddr_axi_s2_o                  : out std_logic_vector(39  downto 0);  -- dahlia_fpga_araddr_axi_s2_i
    fabric_fpga_arburst_axi_s2_o                 : out std_logic_vector(1   downto 0);  -- dahlia_fpga_arburst_axi_s2_i
    fabric_fpga_arcache_axi_s2_o                 : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arcache_axi_s2_i
    fabric_fpga_arid_axi_s2_o                    : out std_logic_vector(11  downto 0);  -- dahlia_fpga_arid_axi_s2_i
    fabric_fpga_arlen_axi_s2_o                   : out std_logic_vector(7   downto 0);  -- dahlia_fpga_arlen_axi_s2_i
    fabric_fpga_arlock_axi_s2_o                  : out std_logic;                       -- dahlia_fpga_arlock_axi_s2_i
    fabric_fpga_arprot_axi_s2_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_arprot_axi_s2_i
    fabric_fpga_arqos_axi_s2_o                   : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arqos_axi_s2_i
    fabric_fpga_arregion_axi_s2_o                : out std_logic_vector(3   downto 0);  -- dahlia_fpga_arregion_axi_s2_i
    fabric_fpga_arsize_axi_s2_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_arsize_axi_s2_i
    fabric_fpga_arvalid_axi_s2_o                 : out std_logic;                       -- dahlia_fpga_arvalid_axi_s2_i
    fabric_fpga_awaddr_axi_s2_o                  : out std_logic_vector(39  downto 0);  -- dahlia_fpga_awaddr_axi_s2_i
    fabric_fpga_awburst_axi_s2_o                 : out std_logic_vector(1   downto 0);  -- dahlia_fpga_awburst_axi_s2_i
    fabric_fpga_awcache_axi_s2_o                 : out std_logic_vector(3   downto 0);  -- dahlia_fpga_awcache_axi_s2_i
    fabric_fpga_awid_axi_s2_o                    : out std_logic_vector(11  downto 0);  -- dahlia_fpga_awid_axi_s2_i
    fabric_fpga_awlen_axi_s2_o                   : out std_logic_vector(7   downto 0);  -- dahlia_fpga_awlen_axi_s2_i
    fabric_fpga_awlock_axi_s2_o                  : out std_logic;                       -- dahlia_fpga_awlock_axi_s2_i
    fabric_fpga_awprot_axi_s2_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_awprot_axi_s2_i
    fabric_fpga_awqos_axi_s2_o                   : out std_logic_vector(3   downto 0);  -- dahlia_fpga_awqos_axi_s2_i
    fabric_fpga_awregion_axi_s2_o                : out std_logic_vector(3   downto 0);  -- dahlia_fpga_awregion_axi_s2_i
    fabric_fpga_awsize_axi_s2_o                  : out std_logic_vector(2   downto 0);  -- dahlia_fpga_awsize_axi_s2_i
    fabric_fpga_bready_axi_s2_o                  : out std_logic;                       -- dahlia_fpga_bready_axi_s2_i
    fabric_fpga_rready_axi_s2_o                  : out std_logic;                       -- dahlia_fpga_rready_axi_s2_i
    fabric_fpga_wdata_axi_s2_o                   : out std_logic_vector(127 downto 0);  -- dahlia_fpga_wdata_axi_s2_i
    fabric_fpga_wlast_axi_s2_o                   : out std_logic;                       -- dahlia_fpga_wlast_axi_s2_i
    fabric_fpga_wstrb_axi_s2_o                   : out std_logic_vector(15  downto 0);  -- dahlia_fpga_wstrb_axi_s2_i
    fabric_fpga_wvalid_axi_s2_o                  : out std_logic;                       -- dahlia_fpga_wvalid_axi_s2_i
    fabric_fpga_awvalid_axi_s2_o                 : out std_logic;                       -- dahlia_fpga_awvalid_axi_s2_i
    fabric_fpga_arready_axi_s2_i                 : in  std_logic;                       -- dahlia_fpga_arready_axi_s2_o
    fabric_fpga_awready_axi_s2_i                 : in  std_logic;                       -- dahlia_fpga_awready_axi_s2_o
    fabric_fpga_bid_axi_s2_i                     : in  std_logic_vector(11  downto 0);  -- dahlia_fpga_bid_axi_s2_o
    fabric_fpga_bresp_axi_s2_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_bresp_axi_s2_o
    fabric_fpga_bvalid_axi_s2_i                  : in  std_logic;                       -- dahlia_fpga_bvalid_axi_s2_o
    fabric_fpga_rdata_axi_s2_i                   : in  std_logic_vector(127 downto 0);  -- dahlia_fpga_rdata_axi_s2_o
    fabric_fpga_rid_axi_s2_i                     : in  std_logic_vector(11  downto 0);  -- dahlia_fpga_rid_axi_s2_o
    fabric_fpga_rlast_axi_s2_i                   : in  std_logic;                       -- dahlia_fpga_rlast_axi_s2_o
    fabric_fpga_rresp_axi_s2_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_rresp_axi_s2_o
    fabric_fpga_rvalid_axi_s2_i                  : in  std_logic;                       -- dahlia_fpga_rvalid_axi_s2_o
    fabric_fpga_wready_axi_s2_i                  : in  std_logic;                       -- dahlia_fpga_wready_axi_s2_o
    fabric_fpga_arready_axi_m1_o                 : out std_logic;                       -- dahlia_fpga_arready_axi_m1_i
    fabric_fpga_awready_axi_m1_o                 : out std_logic;                       -- dahlia_fpga_awready_axi_m1_i
    fabric_fpga_bid_axi_m1_o                     : out std_logic_vector(4   downto 0);  -- dahlia_fpga_bid_axi_m1_i
    fabric_fpga_bresp_axi_m1_o                   : out std_logic_vector(1   downto 0);  -- dahlia_fpga_bresp_axi_m1_i
    fabric_fpga_bvalid_axi_m1_o                  : out std_logic;                       -- dahlia_fpga_bvalid_axi_m1_i
    fabric_fpga_dma_ack_m1_o                     : out std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_ack_m1_i
    fabric_fpga_dma_finish_m1_o                  : out std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_finish_m1_i
    fabric_fpga_rdata_axi_m1_o                   : out std_logic_vector(127 downto 0);  -- dahlia_fpga_rdata_axi_m1_i
    fabric_fpga_rid_axi_m1_o                     : out std_logic_vector(4   downto 0);  -- dahlia_fpga_rid_axi_m1_i
    fabric_fpga_rlast_axi_m1_o                   : out std_logic;                       -- dahlia_fpga_rlast_axi_m1_i
    fabric_fpga_rresp_axi_m1_o                   : out std_logic_vector(1   downto 0);  -- dahlia_fpga_rresp_axi_m1_i
    fabric_fpga_rvalid_axi_m1_o                  : out std_logic;                       -- dahlia_fpga_rvalid_axi_m1_i
    fabric_fpga_wready_axi_m1_o                  : out std_logic;                       -- dahlia_fpga_wready_axi_m1_i
    fabric_fpga_araddr_axi_m1_i                  : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_araddr_axi_m1_o
    fabric_fpga_arburst_axi_m1_i                 : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_arburst_axi_m1_o
    fabric_fpga_arcache_axi_m1_i                 : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_arcache_axi_m1_o
    fabric_fpga_arid_axi_m1_i                    : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_arid_axi_m1_o
    fabric_fpga_arlen_axi_m1_i                   : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_arlen_axi_m1_o
    fabric_fpga_arlock_axi_m1_i                  : in  std_logic;                       -- dahlia_fpga_arlock_axi_m1_o
    fabric_fpga_arprot_axi_m1_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_arprot_axi_m1_o
    fabric_fpga_arqos_axi_m1_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_arqos_axi_m1_o
    fabric_fpga_arsize_axi_m1_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_arsize_axi_m1_o
    fabric_fpga_arvalid_axi_m1_i                 : in  std_logic;                       -- dahlia_fpga_arvalid_axi_m1_o
    fabric_fpga_awaddr_axi_m1_i                  : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_awaddr_axi_m1_o
    fabric_fpga_awburst_axi_m1_i                 : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_awburst_axi_m1_o
    fabric_fpga_awcache_axi_m1_i                 : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_awcache_axi_m1_o
    fabric_fpga_awid_axi_m1_i                    : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_awid_axi_m1_o
    fabric_fpga_awlen_axi_m1_i                   : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_awlen_axi_m1_o
    fabric_fpga_awlock_axi_m1_i                  : in  std_logic;                       -- dahlia_fpga_awlock_axi_m1_o
    fabric_fpga_awprot_axi_m1_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_awprot_axi_m1_o
    fabric_fpga_awqos_axi_m1_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_awqos_axi_m1_o
    fabric_fpga_awsize_axi_m1_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_awsize_axi_m1_o
    fabric_fpga_awvalid_axi_m1_i                 : in  std_logic;                       -- dahlia_fpga_awvalid_axi_m1_o
    fabric_fpga_bready_axi_m1_i                  : in  std_logic;                       -- dahlia_fpga_bready_axi_m1_o
    fabric_fpga_dma_last_m1_i                    : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_last_m1_o
    fabric_fpga_dma_req_m1_i                     : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_req_m1_o
    fabric_fpga_dma_single_m1_i                  : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_single_m1_o
    fabric_fpga_rready_axi_m1_i                  : in  std_logic;                       -- dahlia_fpga_rready_axi_m1_o
    fabric_fpga_wdata_axi_m1_i                   : in  std_logic_vector(127 downto 0);  -- dahlia_fpga_wdata_axi_m1_o
    fabric_fpga_wlast_axi_m1_i                   : in  std_logic;                       -- dahlia_fpga_wlast_axi_m1_o
    fabric_fpga_wstrb_axi_m1_i                   : in  std_logic_vector(15  downto 0);  -- dahlia_fpga_wstrb_axi_m1_o
    fabric_fpga_wvalid_axi_m1_i                  : in  std_logic;                       -- dahlia_fpga_wvalid_axi_m1_o
    fabric_fpga_arready_axi_m2_o                 : out std_logic;                       -- dahlia_fpga_arready_axi_m2_i
    fabric_fpga_awready_axi_m2_o                 : out std_logic;                       -- dahlia_fpga_awready_axi_m2_i
    fabric_fpga_bid_axi_m2_o                     : out std_logic_vector(4   downto 0);  -- dahlia_fpga_bid_axi_m2_i
    fabric_fpga_bresp_axi_m2_o                   : out std_logic_vector(1   downto 0);  -- dahlia_fpga_bresp_axi_m2_i
    fabric_fpga_bvalid_axi_m2_o                  : out std_logic;                       -- dahlia_fpga_bvalid_axi_m2_i
    fabric_fpga_dma_ack_m2_o                     : out std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_ack_m2_i
    fabric_fpga_dma_finish_m2_o                  : out std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_finish_m2_i
    fabric_fpga_rdata_axi_m2_o                   : out std_logic_vector(127 downto 0);  -- dahlia_fpga_rdata_axi_m2_i
    fabric_fpga_rid_axi_m2_o                     : out std_logic_vector(4   downto 0);  -- dahlia_fpga_rid_axi_m2_i
    fabric_fpga_rlast_axi_m2_o                   : out std_logic;                       -- dahlia_fpga_rlast_axi_m2_i
    fabric_fpga_rresp_axi_m2_o                   : out std_logic_vector(1   downto 0);  -- dahlia_fpga_rresp_axi_m2_i
    fabric_fpga_rvalid_axi_m2_o                  : out std_logic;                       -- dahlia_fpga_rvalid_axi_m2_i
    fabric_fpga_wready_axi_m2_o                  : out std_logic;                       -- dahlia_fpga_wready_axi_m2_i
    fabric_fpga_araddr_axi_m2_i                  : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_araddr_axi_m2_o
    fabric_fpga_arburst_axi_m2_i                 : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_arburst_axi_m2_o
    fabric_fpga_arcache_axi_m2_i                 : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_arcache_axi_m2_o
    fabric_fpga_arid_axi_m2_i                    : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_arid_axi_m2_o
    fabric_fpga_arlen_axi_m2_i                   : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_arlen_axi_m2_o
    fabric_fpga_arlock_axi_m2_i                  : in  std_logic;                       -- dahlia_fpga_arlock_axi_m2_o
    fabric_fpga_arprot_axi_m2_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_arprot_axi_m2_o
    fabric_fpga_arqos_axi_m2_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_arqos_axi_m2_o
    fabric_fpga_arsize_axi_m2_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_arsize_axi_m2_o
    fabric_fpga_arvalid_axi_m2_i                 : in  std_logic;                       -- dahlia_fpga_arvalid_axi_m2_o
    fabric_fpga_awaddr_axi_m2_i                  : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_awaddr_axi_m2_o
    fabric_fpga_awburst_axi_m2_i                 : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_awburst_axi_m2_o
    fabric_fpga_awcache_axi_m2_i                 : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_awcache_axi_m2_o
    fabric_fpga_awid_axi_m2_i                    : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_awid_axi_m2_o
    fabric_fpga_awlen_axi_m2_i                   : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_awlen_axi_m2_o
    fabric_fpga_awlock_axi_m2_i                  : in  std_logic;                       -- dahlia_fpga_awlock_axi_m2_o
    fabric_fpga_awprot_axi_m2_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_awprot_axi_m2_o
    fabric_fpga_awqos_axi_m2_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_awqos_axi_m2_o
    fabric_fpga_awsize_axi_m2_i                  : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_awsize_axi_m2_o
    fabric_fpga_awvalid_axi_m2_i                 : in  std_logic;                       -- dahlia_fpga_awvalid_axi_m2_o
    fabric_fpga_bready_axi_m2_i                  : in  std_logic;                       -- dahlia_fpga_bready_axi_m2_o
    fabric_fpga_dma_last_m2_i                    : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_last_m2_o
    fabric_fpga_dma_req_m2_i                     : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_req_m2_o
    fabric_fpga_dma_single_m2_i                  : in  std_logic_vector(5   downto 0);  -- dahlia_fpga_dma_single_m2_o
    fabric_fpga_rready_axi_m2_i                  : in  std_logic;                       -- dahlia_fpga_rready_axi_m2_o
    fabric_fpga_wdata_axi_m2_i                   : in  std_logic_vector(127 downto 0);  -- dahlia_fpga_wdata_axi_m2_o
    fabric_fpga_wlast_axi_m2_i                   : in  std_logic;                       -- dahlia_fpga_wlast_axi_m2_o
    fabric_fpga_wstrb_axi_m2_i                   : in  std_logic_vector(15  downto 0);  -- dahlia_fpga_wstrb_axi_m2_o
    fabric_fpga_wvalid_axi_m2_i                  : in  std_logic;                       -- dahlia_fpga_wvalid_axi_m2_o
    fabric_fpga_ddr0_arready_o                   : out std_logic;                       -- dahlia_fpga_ddr0_arready_i
    fabric_fpga_ddr0_awready_o                   : out std_logic;                       -- dahlia_fpga_ddr0_awready_i
    fabric_fpga_ddr0_bid_o                       : out std_logic_vector(4   downto 0);  -- dahlia_fpga_ddr0_bid_i
    fabric_fpga_ddr0_bresp_o                     : out std_logic_vector(1   downto 0);  -- dahlia_fpga_ddr0_bresp_i
    fabric_fpga_ddr0_bvalid_o                    : out std_logic;                       -- dahlia_fpga_ddr0_bvalid_i
    fabric_fpga_ddr0_rdata_o                     : out std_logic_vector(127 downto 0);  -- dahlia_fpga_ddr0_rdata_i
    fabric_fpga_ddr0_rid_o                       : out std_logic_vector(4   downto 0);  -- dahlia_fpga_ddr0_rid_i
    fabric_fpga_ddr0_rlast_o                     : out std_logic;                       -- dahlia_fpga_ddr0_rlast_i
    fabric_fpga_ddr0_rresp_o                     : out std_logic_vector(1   downto 0);  -- dahlia_fpga_ddr0_rresp_i
    fabric_fpga_ddr0_rvalid_o                    : out std_logic;                       -- dahlia_fpga_ddr0_rvalid_i
    fabric_fpga_ddr0_wready_o                    : out std_logic;                       -- dahlia_fpga_ddr0_wready_i
    fabric_fpga_ddr0_araddr_i                    : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_ddr0_araddr_o
    fabric_fpga_ddr0_arburst_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_ddr0_arburst_o
    fabric_fpga_ddr0_arcache_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_ddr0_arcache_o
    fabric_fpga_ddr0_arid_i                      : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_ddr0_arid_o
    fabric_fpga_ddr0_arlen_i                     : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_ddr0_arlen_o
    fabric_fpga_ddr0_arlock_i                    : in  std_logic;                       -- dahlia_fpga_ddr0_arlock_o
    fabric_fpga_ddr0_arprot_i                    : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_ddr0_arprot_o
    fabric_fpga_ddr0_arqos_i                     : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_ddr0_arqos_o
    fabric_fpga_ddr0_arsize_i                    : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_ddr0_arsize_o
    fabric_fpga_ddr0_arvalid_i                   : in  std_logic;                       -- dahlia_fpga_ddr0_arvalid_o
    fabric_fpga_ddr0_awaddr_i                    : in  std_logic_vector(39  downto 0);  -- dahlia_fpga_ddr0_awaddr_o
    fabric_fpga_ddr0_awburst_i                   : in  std_logic_vector(1   downto 0);  -- dahlia_fpga_ddr0_awburst_o
    fabric_fpga_ddr0_awcache_i                   : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_ddr0_awcache_o
    fabric_fpga_ddr0_awid_i                      : in  std_logic_vector(4   downto 0);  -- dahlia_fpga_ddr0_awid_o
    fabric_fpga_ddr0_awlen_i                     : in  std_logic_vector(7   downto 0);  -- dahlia_fpga_ddr0_awlen_o
    fabric_fpga_ddr0_awlock_i                    : in  std_logic;                       -- dahlia_fpga_ddr0_awlock_o
    fabric_fpga_ddr0_awprot_i                    : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_ddr0_awprot_o
    fabric_fpga_ddr0_awqos_i                     : in  std_logic_vector(3   downto 0);  -- dahlia_fpga_ddr0_awqos_o
    fabric_fpga_ddr0_awsize_i                    : in  std_logic_vector(2   downto 0);  -- dahlia_fpga_ddr0_awsize_o
    fabric_fpga_ddr0_awvalid_i                   : in  std_logic;                       -- dahlia_fpga_ddr0_awvalid_o
    fabric_fpga_ddr0_bready_i                    : in  std_logic;                       -- dahlia_fpga_ddr0_bready_o
    fabric_fpga_ddr0_rready_i                    : in  std_logic;                       -- dahlia_fpga_ddr0_rready_o
    fabric_fpga_ddr0_wdata_i                     : in  std_logic_vector(127 downto 0);  -- dahlia_fpga_ddr0_wdata_o
    fabric_fpga_ddr0_wlast_i                     : in  std_logic;                       -- dahlia_fpga_ddr0_wlast_o
    fabric_fpga_ddr0_wstrb_i                     : in  std_logic_vector(15  downto 0);  -- dahlia_fpga_ddr0_wstrb_o
    fabric_fpga_ddr0_wvalid_i                    : in  std_logic;                       -- dahlia_fpga_ddr0_wvalid_o
    fabric_fpga_paddr_apb_o                      : out std_logic_vector(31  downto 0);  -- dahlia_fpga_paddr_apb_i
    fabric_fpga_penable_apb_o                    : out std_logic;                       -- dahlia_fpga_penable_apb_i
    fabric_fpga_psel_apb_o                       : out std_logic;                       -- dahlia_fpga_psel_apb_i
    fabric_fpga_pwdata_apb_o                     : out std_logic_vector(31  downto 0);  -- dahlia_fpga_pwdata_apb_i
    fabric_fpga_pwrite_apb_o                     : out std_logic;                       -- dahlia_fpga_pwrite_apb_i
    fabric_fpga_prdata_apb_i                     : in  std_logic_vector(31  downto 0);  -- dahlia_fpga_prdata_apb_o
    fabric_fpga_pready_apb_i                     : in  std_logic;                       -- dahlia_fpga_pready_apb_o
    fabric_fpga_pslverr_apb_i                    : in  std_logic;                       -- dahlia_fpga_pslverr_apb_o
    fabric_llpp0_araddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp0_araddr_s_i
    fabric_llpp0_arburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp0_arburst_s_i
    fabric_llpp0_arcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp0_arcache_s_i
    fabric_llpp0_arid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp0_arid_s_i
    fabric_llpp0_arlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp0_arlen_s_i
    fabric_llpp0_arlock_s_o                      : out std_logic;                       -- dahlia_llpp0_arlock_s_i
    fabric_llpp0_arprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp0_arprot_s_i
    fabric_llpp0_arqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp0_arqos_s_i
    fabric_llpp0_arsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp0_arsize_s_i
    fabric_llpp0_arvalid_s_o                     : out std_logic;                       -- dahlia_llpp0_arvalid_s_i
    fabric_llpp0_awaddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp0_awaddr_s_i
    fabric_llpp0_awburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp0_awburst_s_i
    fabric_llpp0_awcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp0_awcache_s_i
    fabric_llpp0_awid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp0_awid_s_i
    fabric_llpp0_awlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp0_awlen_s_i
    fabric_llpp0_awlock_s_o                      : out std_logic;                       -- dahlia_llpp0_awlock_s_i
    fabric_llpp0_awprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp0_awprot_s_i
    fabric_llpp0_awqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp0_awqos_s_i
    fabric_llpp0_awsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp0_awsize_s_i
    fabric_llpp0_awvalid_s_o                     : out std_logic;                       -- dahlia_llpp0_awvalid_s_i
    fabric_llpp0_bready_s_o                      : out std_logic;                       -- dahlia_llpp0_bready_s_i
    fabric_llpp0_rready_s_o                      : out std_logic;                       -- dahlia_llpp0_rready_s_i
    fabric_llpp0_wdata_s_o                       : out std_logic_vector(31  downto 0);  -- dahlia_llpp0_wdata_s_i
    fabric_llpp0_wlast_s_o                       : out std_logic;                       -- dahlia_llpp0_wlast_s_i
    fabric_llpp0_wstrb_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp0_wstrb_s_i
    fabric_llpp0_wvalid_s_o                      : out std_logic;                       -- dahlia_llpp0_wvalid_s_i
    fabric_llpp0_arready_s_i                     : in  std_logic;                       -- dahlia_llpp0_arready_s_o
    fabric_llpp0_awready_s_i                     : in  std_logic;                       -- dahlia_llpp0_awready_s_o
    fabric_llpp0_bid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp0_bid_s_o
    fabric_llpp0_bresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp0_bresp_s_o
    fabric_llpp0_bvalid_s_i                      : in  std_logic;                       -- dahlia_llpp0_bvalid_s_o
    fabric_llpp0_rdata_s_i                       : in  std_logic_vector(31  downto 0);  -- dahlia_llpp0_rdata_s_o
    fabric_llpp0_rid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp0_rid_s_o
    fabric_llpp0_rlast_s_i                       : in  std_logic;                       -- dahlia_llpp0_rlast_s_o
    fabric_llpp0_rresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp0_rresp_s_o
    fabric_llpp0_rvalid_s_i                      : in  std_logic;                       -- dahlia_llpp0_rvalid_s_o
    fabric_llpp0_wready_s_i                      : in  std_logic;                       -- dahlia_llpp0_wready_s_o
    fabric_llpp1_araddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp1_araddr_s_i
    fabric_llpp1_arburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp1_arburst_s_i
    fabric_llpp1_arcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp1_arcache_s_i
    fabric_llpp1_arid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp1_arid_s_i
    fabric_llpp1_arlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp1_arlen_s_i
    fabric_llpp1_arlock_s_o                      : out std_logic;                       -- dahlia_llpp1_arlock_s_i
    fabric_llpp1_arprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp1_arprot_s_i
    fabric_llpp1_arqos_s1_o                      : out std_logic_vector(3   downto 0);  -- dahlia_llpp1_arqos_s1_i
    fabric_llpp1_arsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp1_arsize_s_i
    fabric_llpp1_arvalid_s_o                     : out std_logic;                       -- dahlia_llpp1_arvalid_s_i
    fabric_llpp1_awaddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp1_awaddr_s_i
    fabric_llpp1_awburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp1_awburst_s_i
    fabric_llpp1_awcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp1_awcache_s_i
    fabric_llpp1_awid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp1_awid_s_i
    fabric_llpp1_awlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp1_awlen_s_i
    fabric_llpp1_awlock_s_o                      : out std_logic;                       -- dahlia_llpp1_awlock_s_i
    fabric_llpp1_awprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp1_awprot_s_i
    fabric_llpp1_awqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp1_awqos_s_i
    fabric_llpp1_awsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp1_awsize_s_i
    fabric_llpp1_awvalid_s_o                     : out std_logic;                       -- dahlia_llpp1_awvalid_s_i
    fabric_llpp1_bready_s_o                      : out std_logic;                       -- dahlia_llpp1_bready_s_i
    fabric_llpp1_rready_s_o                      : out std_logic;                       -- dahlia_llpp1_rready_s_i
    fabric_llpp1_wdata_s_o                       : out std_logic_vector(31  downto 0);  -- dahlia_llpp1_wdata_s_i
    fabric_llpp1_wlast_s_o                       : out std_logic;                       -- dahlia_llpp1_wlast_s_i
    fabric_llpp1_wstrb_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp1_wstrb_s_i
    fabric_llpp1_wvalid_s_o                      : out std_logic;                       -- dahlia_llpp1_wvalid_s_i
    fabric_llpp1_arready_s_i                     : in  std_logic;                       -- dahlia_llpp1_arready_s_o
    fabric_llpp1_awready_s_i                     : in  std_logic;                       -- dahlia_llpp1_awready_s_o
    fabric_llpp1_bid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp1_bid_s_o
    fabric_llpp1_bresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp1_bresp_s_o
    fabric_llpp1_bvalid_s_i                      : in  std_logic;                       -- dahlia_llpp1_bvalid_s_o
    fabric_llpp1_rdata_s_i                       : in  std_logic_vector(31  downto 0);  -- dahlia_llpp1_rdata_s_o
    fabric_llpp1_rid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp1_rid_s_o
    fabric_llpp1_rlast_s_i                       : in  std_logic;                       -- dahlia_llpp1_rlast_s_o
    fabric_llpp1_rresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp1_rresp_s_o
    fabric_llpp1_rvalid_s_i                      : in  std_logic;                       -- dahlia_llpp1_rvalid_s_o
    fabric_llpp1_wready_s_i                      : in  std_logic;                       -- dahlia_llpp1_wready_s_o
    fabric_llpp2_araddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp2_araddr_s_i
    fabric_llpp2_arburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp2_arburst_s_i
    fabric_llpp2_arcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp2_arcache_s_i
    fabric_llpp2_arid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp2_arid_s_i
    fabric_llpp2_arlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp2_arlen_s_i
    fabric_llpp2_arlock_s_o                      : out std_logic;                       -- dahlia_llpp2_arlock_s_i
    fabric_llpp2_arprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp2_arprot_s_i
    fabric_llpp2_arqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp2_arqos_s_i
    fabric_llpp2_arsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp2_arsize_s_i
    fabric_llpp2_arvalid_s_o                     : out std_logic;                       -- dahlia_llpp2_arvalid_s_i
    fabric_llpp2_awaddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp2_awaddr_s_i
    fabric_llpp2_awburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp2_awburst_s_i
    fabric_llpp2_awcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp2_awcache_s_i
    fabric_llpp2_awid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp2_awid_s_i
    fabric_llpp2_awlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp2_awlen_s_i
    fabric_llpp2_awlock_s_o                      : out std_logic;                       -- dahlia_llpp2_awlock_s_i
    fabric_llpp2_awprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp2_awprot_s_i
    fabric_llpp2_awqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp2_awqos_s_i
    fabric_llpp2_awsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp2_awsize_s_i
    fabric_llpp2_awvalid_s_o                     : out std_logic;                       -- dahlia_llpp2_awvalid_s_i
    fabric_llpp2_bready_s_o                      : out std_logic;                       -- dahlia_llpp2_bready_s_i
    fabric_llpp2_rready_s_o                      : out std_logic;                       -- dahlia_llpp2_rready_s_i
    fabric_llpp2_wdata_s_o                       : out std_logic_vector(31  downto 0);  -- dahlia_llpp2_wdata_s_i
    fabric_llpp2_wlast_s_o                       : out std_logic;                        -- dahlia_llpp2_wlast_s_i
    fabric_llpp2_wstrb_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp2_wstrb_s_i
    fabric_llpp2_wvalid_s_o                      : out std_logic;                       -- dahlia_llpp2_wvalid_s_i
    fabric_llpp2_arready_s_i                     : in  std_logic;                       -- dahlia_llpp2_arready_s_o
    fabric_llpp2_awready_s_i                     : in  std_logic;                       -- dahlia_llpp2_awready_s_o
    fabric_llpp2_bid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp2_bid_s_o
    fabric_llpp2_bresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp2_bresp_s_o
    fabric_llpp2_bvalid_s_i                      : in  std_logic;                       -- dahlia_llpp2_bvalid_s_o
    fabric_llpp2_rdata_s_i                       : in  std_logic_vector(31  downto 0);  -- dahlia_llpp2_rdata_s_o
    fabric_llpp2_rid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp2_rid_s_o
    fabric_llpp2_rlast_s_i                       : in  std_logic;                       -- dahlia_llpp2_rlast_s_o
    fabric_llpp2_rresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp2_rresp_s_o
    fabric_llpp2_rvalid_s_i                      : in  std_logic;                       -- dahlia_llpp2_rvalid_s_o
    fabric_llpp2_wready_s_i                      : in  std_logic;                       -- dahlia_llpp2_wready_s_o
    fabric_llpp3_araddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp3_araddr_s_i
    fabric_llpp3_arburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp3_arburst_s_i
    fabric_llpp3_arcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp3_arcache_s_i
    fabric_llpp3_arid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp3_arid_s_i
    fabric_llpp3_arlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp3_arlen_s_i
    fabric_llpp3_arlock_s_o                      : out std_logic;                       -- dahlia_llpp3_arlock_s_i
    fabric_llpp3_arprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp3_arprot_s_i
    fabric_llpp3_arqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp3_arqos_s_i
    fabric_llpp3_arsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp3_arsize_s_i
    fabric_llpp3_arvalid_s_o                     : out std_logic;                       -- dahlia_llpp3_arvalid_s_i
    fabric_llpp3_awaddr_s_o                      : out std_logic_vector(31  downto 0);  -- dahlia_llpp3_awaddr_s_i
    fabric_llpp3_awburst_s_o                     : out std_logic_vector(1   downto 0);  -- dahlia_llpp3_awburst_s_i
    fabric_llpp3_awcache_s_o                     : out std_logic_vector(3   downto 0);  -- dahlia_llpp3_awcache_s_i
    fabric_llpp3_awid_s_o                        : out std_logic_vector(11  downto 0);  -- dahlia_llpp3_awid_s_i
    fabric_llpp3_awlen_s_o                       : out std_logic_vector(7   downto 0);  -- dahlia_llpp3_awlen_s_i
    fabric_llpp3_awlock_s_o                      : out std_logic;                       -- dahlia_llpp3_awlock_s_i
    fabric_llpp3_awprot_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp3_awprot_s_i
    fabric_llpp3_awqos_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp3_awqos_s_i
    fabric_llpp3_awsize_s_o                      : out std_logic_vector(2   downto 0);  -- dahlia_llpp3_awsize_s_i
    fabric_llpp3_awvalid_s_o                     : out std_logic;                       -- dahlia_llpp3_awvalid_s_i
    fabric_llpp3_bready_s_o                      : out std_logic;                       -- dahlia_llpp3_bready_s_i
    fabric_llpp3_rready_s_o                      : out std_logic;                       -- dahlia_llpp3_rready_s_i
    fabric_llpp3_wdata_s_o                       : out std_logic_vector(31  downto 0);  -- dahlia_llpp3_wdata_s_i
    fabric_llpp3_wlast_s_o                       : out std_logic;                       -- dahlia_llpp3_wlast_s_i
    fabric_llpp3_wstrb_s_o                       : out std_logic_vector(3   downto 0);  -- dahlia_llpp3_wstrb_s_i
    fabric_llpp3_wvalid_s_o                      : out std_logic;                       -- dahlia_llpp3_wvalid_s_i
    fabric_llpp3_arready_s_i                     : in  std_logic;                       -- dahlia_llpp3_arready_s_o
    fabric_llpp3_awready_s_i                     : in  std_logic;                       -- dahlia_llpp3_awready_s_o
    fabric_llpp3_bid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp3_bid_s_o
    fabric_llpp3_bresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp3_bresp_s_o
    fabric_llpp3_bvalid_s_i                      : in  std_logic;                       -- dahlia_llpp3_bvalid_s_o
    fabric_llpp3_rdata_s_i                       : in  std_logic_vector(31  downto 0);  -- dahlia_llpp3_rdata_s_o
    fabric_llpp3_rid_s_i                         : in  std_logic_vector(11  downto 0);  -- dahlia_llpp3_rid_s_o
    fabric_llpp3_rlast_s_i                       : in  std_logic;                       -- dahlia_llpp3_rlast_s_o
    fabric_llpp3_rresp_s_i                       : in  std_logic_vector(1   downto 0);  -- dahlia_llpp3_rresp_s_o
    fabric_llpp3_rvalid_s_i                      : in  std_logic;                       -- dahlia_llpp3_rvalid_s_o
    fabric_llpp3_wready_s_i                      : in  std_logic;                       -- dahlia_llpp3_wready_s_o
    fabric_qos_pprdata_o                         : out std_logic_vector(31  downto 0);  -- dahlia_qos_pprdata_i
    fabric_qos_ppready_o                         : out std_logic;                       -- dahlia_qos_ppready_i
    fabric_qos_ppslverr_o                        : out std_logic;                       -- dahlia_qos_ppslverr_i
    fabric_qos_pclk_i                            : in  std_logic;                       -- dahlia_qos_pclk_o
    fabric_qos_ppaddr_i                          : in  std_logic_vector(31  downto 0);  -- dahlia_qos_ppaddr_o
    fabric_qos_ppenable_i                        : in  std_logic;                       -- dahlia_qos_ppenable_o
    fabric_qos_ppwdata_i                         : in  std_logic_vector(31  downto 0);  -- dahlia_qos_ppwdata_o
    fabric_qos_ppwrite_i                         : in  std_logic;                       -- dahlia_qos_ppwrite_o
    fabric_qos_presetn_i                         : in  std_logic;                       -- dahlia_qos_presetn_o
    fabric_qos_psel_i                            : in  std_logic;                       -- dahlia_qos_psel_o
    fabric_tnd_hssl_flushin_o                    : out std_logic;                       -- dahlia_tnd_hssl_flushin_i
    fabric_tnd_hssl_trigin_o                     : out std_logic;                       -- dahlia_tnd_hssl_trigin_i
    fabric_tnd_fpga_apb_master_paddr_o           : out std_logic_vector(31  downto 0);  -- dahlia_tnd_fpga_apb_master_paddr_i
    fabric_tnd_fpga_apb_master_penable_o         : out std_logic;                       -- dahlia_tnd_fpga_apb_master_penable_i
    fabric_tnd_fpga_apb_master_psel_o            : out std_logic;                       -- dahlia_tnd_fpga_apb_master_psel_i
    fabric_tnd_fpga_apb_master_pwdata_o          : out std_logic_vector(31  downto 0);  -- dahlia_tnd_fpga_apb_master_pwdata_i
    fabric_tnd_fpga_apb_master_pwrite_o          : out std_logic;                       -- dahlia_tnd_fpga_apb_master_pwrite_i
    fabric_tnd_fpga_atb_master_afvalid_o         : out std_logic;                       -- dahlia_tnd_fpga_atb_master_afvalid_i
    fabric_tnd_fpga_atb_master_atready_o         : out std_logic;                       -- dahlia_tnd_fpga_atb_master_atready_i
    fabric_tnd_fpga_atb_master_syncreq_o         : out std_logic;                       -- dahlia_tnd_fpga_atb_master_syncreq_i
    fabric_tnd_hssl_apb_master_paddr_o           : out std_logic_vector(31  downto 0);  -- dahlia_tnd_hssl_apb_master_paddr_i
    fabric_tnd_hssl_apb_master_penable_o         : out std_logic;                       -- dahlia_tnd_hssl_apb_master_penable_i
    fabric_tnd_hssl_apb_master_psel_o            : out std_logic;                       -- dahlia_tnd_hssl_apb_master_psel_i
    fabric_tnd_hssl_apb_master_pwdata_o          : out std_logic_vector(31  downto 0);  -- dahlia_tnd_hssl_apb_master_pwdata_i
    fabric_tnd_hssl_apb_master_pwrite_o          : out std_logic;                       -- dahlia_tnd_hssl_apb_master_pwrite_i
    fabric_tnd_hssl_atb_master_afready_o         : out std_logic;                       -- dahlia_tnd_hssl_atb_master_afready_i
    fabric_tnd_hssl_atb_master_atbytes_o         : out std_logic_vector(3   downto 0);  -- dahlia_tnd_hssl_atb_master_atbytes_i
    fabric_tnd_hssl_atb_master_atdata_o          : out std_logic_vector(127 downto 0);  -- dahlia_tnd_hssl_atb_master_atdata_i
    fabric_tnd_hssl_atb_master_atid_o            : out std_logic_vector(6   downto 0);  -- dahlia_tnd_hssl_atb_master_atid_i
    fabric_tnd_hssl_atb_master_atvalid_o         : out std_logic;                       -- dahlia_tnd_hssl_atb_master_atvalid_i
    fabric_tnd_trace_clk_traceoutportintf_o      : out std_logic;                       -- dahlia_tnd_trace_clk_traceoutportintf_i
    fabric_tnd_trace_ctl_traceoutportintf_o      : out std_logic;                       -- dahlia_tnd_trace_ctl_traceoutportintf_i
    fabric_tnd_trace_data_traceoutportintf_o     : out std_logic_vector(31  downto 0);  -- dahlia_tnd_trace_data_traceoutportintf_i
    fabric_tsvalue_tsgen_fpga_o                  : out std_logic_vector(63  downto 0);  -- dahlia_tsvalue_tsgen_fpga_i
    fabric_tnd_fpga_apb_master_prdata_i          : in  std_logic_vector(31  downto 0);  -- dahlia_tnd_fpga_apb_master_prdata_o
    fabric_tnd_fpga_apb_master_pready_i          : in  std_logic;                       -- dahlia_tnd_fpga_apb_master_pready_o
    fabric_tnd_fpga_apb_master_pslverr_i         : in  std_logic;                       -- dahlia_tnd_fpga_apb_master_pslverr_o
    fabric_tnd_fpga_atb_master_afready_i         : in  std_logic;                       -- dahlia_tnd_fpga_atb_master_afready_o
    fabric_tnd_fpga_atb_master_atbytes_i         : in  std_logic_vector(3   downto 0);  -- dahlia_tnd_fpga_atb_master_atbytes_o
    fabric_tnd_fpga_atb_master_atdata_i          : in  std_logic_vector(127 downto 0);  -- dahlia_tnd_fpga_atb_master_atdata_o
    fabric_tnd_fpga_atb_master_atid_i            : in  std_logic_vector(6   downto 0);  -- dahlia_tnd_fpga_atb_master_atid_o
    fabric_tnd_fpga_atb_master_atvalid_i         : in  std_logic;                       -- dahlia_tnd_fpga_atb_master_atvalid_o
    fabric_tnd_hssl_apb_master_prdata_i          : in  std_logic_vector(31  downto 0);  -- dahlia_tnd_hssl_apb_master_prdata_o
    fabric_tnd_hssl_apb_master_pready_i          : in  std_logic;                       -- dahlia_tnd_hssl_apb_master_pready_o
    fabric_tnd_hssl_apb_master_pslverr_i         : in  std_logic;                       -- dahlia_tnd_hssl_apb_master_pslverr_o
    fabric_tnd_hssl_atb_master_afvalid_i         : in  std_logic;                       -- dahlia_tnd_hssl_atb_master_afvalid_o
    fabric_tnd_hssl_atb_master_atready_i         : in  std_logic;                       -- dahlia_tnd_hssl_atb_master_atready_o
    fabric_tnd_hssl_atb_master_syncreq_i         : in  std_logic;                       -- dahlia_tnd_hssl_atb_master_syncreq_o
    fabric_watchdog0_signal_0_o                  : out std_logic;                       -- dahlia_watchdog0_signal_0_i
    fabric_watchdog0_signal_1_o                  : out std_logic;                       -- dahlia_watchdog0_signal_1_i
    fabric_watchdog1_signal_0_o                  : out std_logic;                       -- dahlia_watchdog1_signal_0_i
    fabric_watchdog1_signal_1_o                  : out std_logic;                       -- dahlia_watchdog1_signal_1_i
    fabric_watchdog2_signal_0_o                  : out std_logic;                       -- dahlia_watchdog2_signal_0_i
    fabric_watchdog2_signal_1_o                  : out std_logic;                       -- dahlia_watchdog2_signal_1_i
    fabric_watchdog3_signal_0_o                  : out std_logic;                       -- dahlia_watchdog3_signal_0_i
    fabric_watchdog3_signal_1_o                  : out std_logic;                       -- dahlia_watchdog3_signal_1_i
    fabric_tst_pll_lock_o                        : out std_logic_vector(6   downto 0);  -- dahlia_tst_pll_lock_i
    fabric_soc_mon_sensor_alarm_o                : out std_logic;                       -- dahlia_soc_mon_sensor_alarm_i
    fabric_erom_fpga_cpu0_dbgen_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu0_dbgen_o
    fabric_erom_fpga_cpu0_hiden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu0_hiden_o
    fabric_erom_fpga_cpu0_hniden_i               : in  std_logic;                       -- dahlia_erom_fpga_cpu0_hniden_o
    fabric_erom_fpga_cpu0_niden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu0_niden_o
    fabric_erom_fpga_cpu1_dbgen_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu1_dbgen_o
    fabric_erom_fpga_cpu1_hiden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu1_hiden_o
    fabric_erom_fpga_cpu1_hniden_i               : in  std_logic;                       -- dahlia_erom_fpga_cpu1_hniden_o
    fabric_erom_fpga_cpu1_niden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu1_niden_o
    fabric_erom_fpga_cpu2_dbgen_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu2_dbgen_o
    fabric_erom_fpga_cpu2_hiden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu2_hiden_o
    fabric_erom_fpga_cpu2_hniden_i               : in  std_logic;                       -- dahlia_erom_fpga_cpu2_hniden_o
    fabric_erom_fpga_cpu2_niden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu2_niden_o
    fabric_erom_fpga_cpu3_dbgen_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu3_dbgen_o
    fabric_erom_fpga_cpu3_hiden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu3_hiden_o
    fabric_erom_fpga_cpu3_hniden_i               : in  std_logic;                       -- dahlia_erom_fpga_cpu3_hniden_o
    fabric_erom_fpga_cpu3_niden_i                : in  std_logic;                       -- dahlia_erom_fpga_cpu3_niden_o
    fabric_erom_fpga_cs_dbgen_i                  : in  std_logic;                       -- dahlia_erom_fpga_cs_dbgen_o
    fabric_erom_fpga_cs_niden_i                  : in  std_logic;                       -- dahlia_erom_fpga_cs_niden_o
    fabric_erom_fpga_cs_deviceen_i               : in  std_logic;                       -- dahlia_erom_fpga_cs_deviceen_o
    fabric_erom_fpga_cs_rst_n_i                  : in  std_logic;                       -- dahlia_erom_fpga_cs_rst_n_o
    fabric_erom_fpga_debug_en_i                  : in  std_logic;                       -- dahlia_erom_fpga_debug_en_o
    fabric_enable_TMR_i                          : in  std_logic_vector(3   downto 0)
);
end NX_SOC_INTERFACE_WRAP;

architecture NX_RTL of NX_SOC_INTERFACE_WRAP is
begin

    inst_NX_SOC : NX_SOC_INTERFACE
    port map (
         fabric_lowskew_o1                           =>  fabric_lowskew_o(0)
       , fabric_lowskew_o2                           =>  fabric_lowskew_o(1)
       , fabric_lowskew_i1                           =>  fabric_lowskew_i(0)
       , fabric_lowskew_i2                           =>  fabric_lowskew_i(1)
       , fabric_lowskew_i3                           =>  fabric_lowskew_i(2)
       , fabric_lowskew_i4                           =>  fabric_lowskew_i(3)
       , fabric_lowskew_i5                           =>  fabric_lowskew_i(4)
       , fabric_lowskew_i6                           =>  fabric_lowskew_i(5)
       , fabric_lowskew_i7                           =>  fabric_lowskew_i(6)
       , fabric_lowskew_i8                           =>  fabric_lowskew_i(7)
       , fabric_lowskew_i9                           =>  fabric_lowskew_i(8)
       , fabric_lowskew_i10                          =>  fabric_lowskew_i(9)
       , fabric_fpga_nic_rstn_i1                     =>  fabric_fpga_nic_rstn_i(0)
       , fabric_fpga_nic_rstn_i2                     =>  fabric_fpga_nic_rstn_i(1)
       , fabric_fpga_nic_rstn_i3                     =>  fabric_fpga_nic_rstn_i(2)
       , fabric_fpga_nic_rstn_i4                     =>  fabric_fpga_nic_rstn_i(3)
       , fabric_fpga_nic_rstn_i5                     =>  fabric_fpga_nic_rstn_i(4)
       , fabric_fpga_nic_rstn_i6                     =>  fabric_fpga_nic_rstn_i(5)
       , fabric_fpga_nic_rstn_i7                     =>  fabric_fpga_nic_rstn_i(6)
       , fabric_fpga_nic_rstn_i8                     =>  fabric_fpga_nic_rstn_i(7)
       , fabric_fpga_nic_rstn_i9                     =>  fabric_fpga_nic_rstn_i(8)
       , fabric_fpga_nic_rstn_i10                    =>  fabric_fpga_nic_rstn_i(9)
       , fabric_fpga_pmrstn_i                        =>  fabric_fpga_pmrstn_i
       , fabric_fpga_sysrstn_i                       =>  fabric_fpga_sysrstn_i
       , fabric_fpga_trigger_in_o1                   =>  fabric_fpga_trigger_in_o(0)
       , fabric_fpga_trigger_in_o2                   =>  fabric_fpga_trigger_in_o(1)
       , fabric_fpga_trigger_in_o3                   =>  fabric_fpga_trigger_in_o(2)
       , fabric_fpga_trigger_in_o4                   =>  fabric_fpga_trigger_in_o(3)
       , fabric_fpga_trigger_in_o5                   =>  fabric_fpga_trigger_in_o(4)
       , fabric_fpga_trigger_in_o6                   =>  fabric_fpga_trigger_in_o(5)
       , fabric_fpga_trigger_in_o7                   =>  fabric_fpga_trigger_in_o(6)
       , fabric_fpga_trigger_in_o8                   =>  fabric_fpga_trigger_in_o(7)
       , fabric_fpga_trigger_out_i1                  =>  fabric_fpga_trigger_out_i(0)
       , fabric_fpga_trigger_out_i2                  =>  fabric_fpga_trigger_out_i(1)
       , fabric_fpga_trigger_out_i3                  =>  fabric_fpga_trigger_out_i(2)
       , fabric_fpga_trigger_out_i4                  =>  fabric_fpga_trigger_out_i(3)
       , fabric_fpga_trigger_out_i5                  =>  fabric_fpga_trigger_out_i(4)
       , fabric_fpga_trigger_out_i6                  =>  fabric_fpga_trigger_out_i(5)
       , fabric_fpga_trigger_out_i7                  =>  fabric_fpga_trigger_out_i(6)
       , fabric_fpga_trigger_out_i8                  =>  fabric_fpga_trigger_out_i(7)
       , fabric_fpga_interrupt_in_i1                 =>  fabric_fpga_interrupt_in_i(0)
       , fabric_fpga_interrupt_in_i2                 =>  fabric_fpga_interrupt_in_i(1)
       , fabric_fpga_interrupt_in_i3                 =>  fabric_fpga_interrupt_in_i(2)
       , fabric_fpga_interrupt_in_i4                 =>  fabric_fpga_interrupt_in_i(3)
       , fabric_fpga_interrupt_in_i5                 =>  fabric_fpga_interrupt_in_i(4)
       , fabric_fpga_interrupt_in_i6                 =>  fabric_fpga_interrupt_in_i(5)
       , fabric_fpga_interrupt_in_i7                 =>  fabric_fpga_interrupt_in_i(6)
       , fabric_fpga_interrupt_in_i8                 =>  fabric_fpga_interrupt_in_i(7)
       , fabric_fpga_interrupt_in_i9                 =>  fabric_fpga_interrupt_in_i(8)
       , fabric_fpga_interrupt_in_i10                =>  fabric_fpga_interrupt_in_i(9)
       , fabric_fpga_interrupt_in_i11                =>  fabric_fpga_interrupt_in_i(10)
       , fabric_fpga_interrupt_in_i12                =>  fabric_fpga_interrupt_in_i(11)
       , fabric_fpga_interrupt_in_i13                =>  fabric_fpga_interrupt_in_i(12)
       , fabric_fpga_interrupt_in_i14                =>  fabric_fpga_interrupt_in_i(13)
       , fabric_fpga_interrupt_in_i15                =>  fabric_fpga_interrupt_in_i(14)
       , fabric_fpga_interrupt_in_i16                =>  fabric_fpga_interrupt_in_i(15)
       , fabric_fpga_interrupt_in_i17                =>  fabric_fpga_interrupt_in_i(16)
       , fabric_fpga_interrupt_in_i18                =>  fabric_fpga_interrupt_in_i(17)
       , fabric_fpga_interrupt_in_i19                =>  fabric_fpga_interrupt_in_i(18)
       , fabric_fpga_interrupt_in_i20                =>  fabric_fpga_interrupt_in_i(19)
       , fabric_fpga_interrupt_in_i21                =>  fabric_fpga_interrupt_in_i(20)
       , fabric_fpga_interrupt_in_i22                =>  fabric_fpga_interrupt_in_i(21)
       , fabric_fpga_interrupt_in_i23                =>  fabric_fpga_interrupt_in_i(22)
       , fabric_fpga_interrupt_in_i24                =>  fabric_fpga_interrupt_in_i(23)
       , fabric_fpga_interrupt_in_i25                =>  fabric_fpga_interrupt_in_i(24)
       , fabric_fpga_interrupt_in_i26                =>  fabric_fpga_interrupt_in_i(25)
       , fabric_fpga_interrupt_in_i27                =>  fabric_fpga_interrupt_in_i(26)
       , fabric_fpga_interrupt_in_i28                =>  fabric_fpga_interrupt_in_i(27)
       , fabric_fpga_interrupt_in_i29                =>  fabric_fpga_interrupt_in_i(28)
       , fabric_fpga_interrupt_in_i30                =>  fabric_fpga_interrupt_in_i(29)
       , fabric_fpga_interrupt_in_i31                =>  fabric_fpga_interrupt_in_i(30)
       , fabric_fpga_interrupt_in_i32                =>  fabric_fpga_interrupt_in_i(31)
       , fabric_fpga_interrupt_in_i33                =>  fabric_fpga_interrupt_in_i(32)
       , fabric_fpga_interrupt_in_i34                =>  fabric_fpga_interrupt_in_i(33)
       , fabric_fpga_interrupt_in_i35                =>  fabric_fpga_interrupt_in_i(34)
       , fabric_fpga_interrupt_in_i36                =>  fabric_fpga_interrupt_in_i(35)
       , fabric_fpga_interrupt_in_i37                =>  fabric_fpga_interrupt_in_i(36)
       , fabric_fpga_interrupt_in_i38                =>  fabric_fpga_interrupt_in_i(37)
       , fabric_fpga_interrupt_in_i39                =>  fabric_fpga_interrupt_in_i(38)
       , fabric_fpga_interrupt_in_i40                =>  fabric_fpga_interrupt_in_i(39)
       , fabric_fpga_interrupt_in_i41                =>  fabric_fpga_interrupt_in_i(40)
       , fabric_fpga_interrupt_in_i42                =>  fabric_fpga_interrupt_in_i(41)
       , fabric_fpga_interrupt_in_i43                =>  fabric_fpga_interrupt_in_i(42)
       , fabric_fpga_interrupt_in_i44                =>  fabric_fpga_interrupt_in_i(43)
       , fabric_fpga_interrupt_in_i45                =>  fabric_fpga_interrupt_in_i(44)
       , fabric_fpga_interrupt_in_i46                =>  fabric_fpga_interrupt_in_i(45)
       , fabric_fpga_interrupt_in_i47                =>  fabric_fpga_interrupt_in_i(46)
       , fabric_fpga_interrupt_in_i48                =>  fabric_fpga_interrupt_in_i(47)
       , fabric_fpga_interrupt_in_i49                =>  fabric_fpga_interrupt_in_i(48)
       , fabric_fpga_interrupt_in_i50                =>  fabric_fpga_interrupt_in_i(49)
       , fabric_fpga_interrupt_in_i51                =>  fabric_fpga_interrupt_in_i(50)
       , fabric_fpga_interrupt_in_i52                =>  fabric_fpga_interrupt_in_i(51)
       , fabric_fpga_interrupt_in_i53                =>  fabric_fpga_interrupt_in_i(52)
       , fabric_fpga_interrupt_in_i54                =>  fabric_fpga_interrupt_in_i(53)
       , fabric_fpga_interrupt_in_i55                =>  fabric_fpga_interrupt_in_i(54)
       , fabric_fpga_interrupt_in_i56                =>  fabric_fpga_interrupt_in_i(55)
       , fabric_fpga_interrupt_in_i57                =>  fabric_fpga_interrupt_in_i(56)
       , fabric_fpga_interrupt_in_i58                =>  fabric_fpga_interrupt_in_i(57)
       , fabric_fpga_interrupt_in_i59                =>  fabric_fpga_interrupt_in_i(58)
       , fabric_fpga_interrupt_in_i60                =>  fabric_fpga_interrupt_in_i(59)
       , fabric_fpga_interrupt_in_i61                =>  fabric_fpga_interrupt_in_i(60)
       , fabric_fpga_interrupt_in_i62                =>  fabric_fpga_interrupt_in_i(61)
       , fabric_fpga_interrupt_in_i63                =>  fabric_fpga_interrupt_in_i(62)
       , fabric_fpga_interrupt_in_i64                =>  fabric_fpga_interrupt_in_i(63)
       , fabric_fpga_interrupt_in_i65                =>  fabric_fpga_interrupt_in_i(64)
       , fabric_fpga_interrupt_in_i66                =>  fabric_fpga_interrupt_in_i(65)
       , fabric_fpga_interrupt_in_i67                =>  fabric_fpga_interrupt_in_i(66)
       , fabric_fpga_interrupt_in_i68                =>  fabric_fpga_interrupt_in_i(67)
       , fabric_fpga_interrupt_in_i69                =>  fabric_fpga_interrupt_in_i(68)
       , fabric_fpga_interrupt_in_i70                =>  fabric_fpga_interrupt_in_i(69)
       , fabric_fpga_interrupt_in_i71                =>  fabric_fpga_interrupt_in_i(70)
       , fabric_fpga_interrupt_in_i72                =>  fabric_fpga_interrupt_in_i(71)
       , fabric_fpga_interrupt_in_i73                =>  fabric_fpga_interrupt_in_i(72)
       , fabric_fpga_interrupt_in_i74                =>  fabric_fpga_interrupt_in_i(73)
       , fabric_fpga_interrupt_in_i75                =>  fabric_fpga_interrupt_in_i(74)
       , fabric_fpga_interrupt_in_i76                =>  fabric_fpga_interrupt_in_i(75)
       , fabric_fpga_interrupt_in_i77                =>  fabric_fpga_interrupt_in_i(76)
       , fabric_fpga_interrupt_in_i78                =>  fabric_fpga_interrupt_in_i(77)
       , fabric_fpga_interrupt_in_i79                =>  fabric_fpga_interrupt_in_i(78)
       , fabric_fpga_interrupt_in_i80                =>  fabric_fpga_interrupt_in_i(79)
       , fabric_fpga_interrupt_in_i81                =>  fabric_fpga_interrupt_in_i(80)
       , fabric_fpga_interrupt_in_i82                =>  fabric_fpga_interrupt_in_i(81)
       , fabric_fpga_interrupt_in_i83                =>  fabric_fpga_interrupt_in_i(82)
       , fabric_fpga_interrupt_in_i84                =>  fabric_fpga_interrupt_in_i(83)
       , fabric_fpga_interrupt_in_i85                =>  fabric_fpga_interrupt_in_i(84)
       , fabric_fpga_interrupt_in_i86                =>  fabric_fpga_interrupt_in_i(85)
       , fabric_fpga_interrupt_in_i87                =>  fabric_fpga_interrupt_in_i(86)
       , fabric_fpga_interrupt_in_i88                =>  fabric_fpga_interrupt_in_i(87)
       , fabric_fpga_interrupt_in_i89                =>  fabric_fpga_interrupt_in_i(88)
       , fabric_fpga_interrupt_in_i90                =>  fabric_fpga_interrupt_in_i(89)
       , fabric_fpga_interrupt_in_i91                =>  fabric_fpga_interrupt_in_i(90)
       , fabric_fpga_interrupt_in_i92                =>  fabric_fpga_interrupt_in_i(91)
       , fabric_fpga_interrupt_in_i93                =>  fabric_fpga_interrupt_in_i(92)
       , fabric_fpga_interrupt_in_i94                =>  fabric_fpga_interrupt_in_i(93)
       , fabric_fpga_interrupt_in_i95                =>  fabric_fpga_interrupt_in_i(94)
       , fabric_fpga_interrupt_in_i96                =>  fabric_fpga_interrupt_in_i(95)
       , fabric_fpga_interrupt_in_i97                =>  fabric_fpga_interrupt_in_i(96)
       , fabric_fpga_interrupt_in_i98                =>  fabric_fpga_interrupt_in_i(97)
       , fabric_fpga_interrupt_in_i99                =>  fabric_fpga_interrupt_in_i(98)
       , fabric_fpga_interrupt_in_i100               =>  fabric_fpga_interrupt_in_i(99)
       , fabric_fpga_interrupt_in_i101               =>  fabric_fpga_interrupt_in_i(100)
       , fabric_fpga_interrupt_in_i102               =>  fabric_fpga_interrupt_in_i(101)
       , fabric_fpga_interrupt_in_i103               =>  fabric_fpga_interrupt_in_i(102)
       , fabric_fpga_interrupt_in_i104               =>  fabric_fpga_interrupt_in_i(103)
       , fabric_fpga_interrupt_in_i105               =>  fabric_fpga_interrupt_in_i(104)
       , fabric_fpga_interrupt_in_i106               =>  fabric_fpga_interrupt_in_i(105)
       , fabric_fpga_interrupt_in_i107               =>  fabric_fpga_interrupt_in_i(106)
       , fabric_fpga_interrupt_in_i108               =>  fabric_fpga_interrupt_in_i(107)
       , fabric_fpga_interrupt_in_i109               =>  fabric_fpga_interrupt_in_i(108)
       , fabric_fpga_interrupt_in_i110               =>  fabric_fpga_interrupt_in_i(109)
       , fabric_fpga_interrupt_in_i111               =>  fabric_fpga_interrupt_in_i(110)
       , fabric_fpga_interrupt_in_i112               =>  fabric_fpga_interrupt_in_i(111)
       , fabric_fpga_interrupt_in_i113               =>  fabric_fpga_interrupt_in_i(112)
       , fabric_fpga_interrupt_in_i114               =>  fabric_fpga_interrupt_in_i(113)
       , fabric_fpga_interrupt_in_i115               =>  fabric_fpga_interrupt_in_i(114)
       , fabric_fpga_interrupt_in_i116               =>  fabric_fpga_interrupt_in_i(115)
       , fabric_fpga_interrupt_in_i117               =>  fabric_fpga_interrupt_in_i(116)
       , fabric_fpga_interrupt_in_i118               =>  fabric_fpga_interrupt_in_i(117)
       , fabric_fpga_interrupt_in_i119               =>  fabric_fpga_interrupt_in_i(118)
       , fabric_fpga_interrupt_in_i120               =>  fabric_fpga_interrupt_in_i(119)
       , fabric_sysc_hold_on_debug_i                 =>  fabric_sysc_hold_on_debug_i
       , fabric_fpga_events60_i1                     =>  fabric_fpga_events60_i(0)
       , fabric_fpga_events60_i2                     =>  fabric_fpga_events60_i(1)
       , fabric_fpga_events60_i3                     =>  fabric_fpga_events60_i(2)
       , fabric_fpga_events60_i4                     =>  fabric_fpga_events60_i(3)
       , fabric_fpga_events60_i5                     =>  fabric_fpga_events60_i(4)
       , fabric_fpga_events60_i6                     =>  fabric_fpga_events60_i(5)
       , fabric_fpga_events60_i7                     =>  fabric_fpga_events60_i(6)
       , fabric_fpga_events60_i8                     =>  fabric_fpga_events60_i(7)
       , fabric_fpga_events60_i9                     =>  fabric_fpga_events60_i(8)
       , fabric_fpga_events60_i10                    =>  fabric_fpga_events60_i(9)
       , fabric_fpga_events60_i11                    =>  fabric_fpga_events60_i(10)
       , fabric_fpga_events60_i12                    =>  fabric_fpga_events60_i(11)
       , fabric_fpga_events60_i13                    =>  fabric_fpga_events60_i(12)
       , fabric_fpga_events60_i14                    =>  fabric_fpga_events60_i(13)
       , fabric_fpga_events60_i15                    =>  fabric_fpga_events60_i(14)
       , fabric_fpga_events60_i16                    =>  fabric_fpga_events60_i(15)
       , fabric_fpga_events60_i17                    =>  fabric_fpga_events60_i(16)
       , fabric_fpga_events60_i18                    =>  fabric_fpga_events60_i(17)
       , fabric_fpga_events60_i19                    =>  fabric_fpga_events60_i(18)
       , fabric_fpga_events60_i20                    =>  fabric_fpga_events60_i(19)
       , fabric_fpga_events60_i21                    =>  fabric_fpga_events60_i(20)
       , fabric_fpga_events60_i22                    =>  fabric_fpga_events60_i(21)
       , fabric_fpga_events60_i23                    =>  fabric_fpga_events60_i(22)
       , fabric_fpga_events60_i24                    =>  fabric_fpga_events60_i(23)
       , fabric_fpga_events60_i25                    =>  fabric_fpga_events60_i(24)
       , fabric_fpga_events60_i26                    =>  fabric_fpga_events60_i(25)
       , fabric_fpga_events60_i27                    =>  fabric_fpga_events60_i(26)
       , fabric_fpga_events60_i28                    =>  fabric_fpga_events60_i(27)
       , fabric_fpga_events60_i29                    =>  fabric_fpga_events60_i(28)
       , fabric_fpga_events60_i30                    =>  fabric_fpga_events60_i(29)
       , fabric_fpga_events60_i31                    =>  fabric_fpga_events60_i(30)
       , fabric_fpga_events60_i32                    =>  fabric_fpga_events60_i(31)
       , fabric_fpga_events60_i33                    =>  fabric_fpga_events60_i(32)
       , fabric_fpga_events60_i34                    =>  fabric_fpga_events60_i(33)
       , fabric_fpga_events60_i35                    =>  fabric_fpga_events60_i(34)
       , fabric_fpga_events60_i36                    =>  fabric_fpga_events60_i(35)
       , fabric_fpga_events60_i37                    =>  fabric_fpga_events60_i(36)
       , fabric_fpga_events60_i38                    =>  fabric_fpga_events60_i(37)
       , fabric_fpga_events60_i39                    =>  fabric_fpga_events60_i(38)
       , fabric_fpga_events60_i40                    =>  fabric_fpga_events60_i(39)
       , fabric_fpga_events60_i41                    =>  fabric_fpga_events60_i(40)
       , fabric_fpga_events60_i42                    =>  fabric_fpga_events60_i(41)
       , fabric_fpga_events60_i43                    =>  fabric_fpga_events60_i(42)
       , fabric_fpga_events60_i44                    =>  fabric_fpga_events60_i(43)
       , fabric_fpga_events60_i45                    =>  fabric_fpga_events60_i(44)
       , fabric_fpga_events60_i46                    =>  fabric_fpga_events60_i(45)
       , fabric_fpga_events60_i47                    =>  fabric_fpga_events60_i(46)
       , fabric_fpga_events60_i48                    =>  fabric_fpga_events60_i(47)
       , fabric_fpga_events60_i49                    =>  fabric_fpga_events60_i(48)
       , fabric_fpga_events60_i50                    =>  fabric_fpga_events60_i(49)
       , fabric_fpga_events60_i51                    =>  fabric_fpga_events60_i(50)
       , fabric_fpga_events60_i52                    =>  fabric_fpga_events60_i(51)
       , fabric_fpga_events60_i53                    =>  fabric_fpga_events60_i(52)
       , fabric_fpga_events60_i54                    =>  fabric_fpga_events60_i(53)
       , fabric_fpga_events60_i55                    =>  fabric_fpga_events60_i(54)
       , fabric_fpga_events60_i56                    =>  fabric_fpga_events60_i(55)
       , fabric_fpga_events60_i57                    =>  fabric_fpga_events60_i(56)
       , fabric_fpga_events60_i58                    =>  fabric_fpga_events60_i(57)
       , fabric_fpga_events60_i59                    =>  fabric_fpga_events60_i(58)
       , fabric_fpga_events60_i60                    =>  fabric_fpga_events60_i(59)
       , fabric_fpga_araddr_axi_s1_o1                =>  fabric_fpga_araddr_axi_s1_o(0)
       , fabric_fpga_araddr_axi_s1_o2                =>  fabric_fpga_araddr_axi_s1_o(1)
       , fabric_fpga_araddr_axi_s1_o3                =>  fabric_fpga_araddr_axi_s1_o(2)
       , fabric_fpga_araddr_axi_s1_o4                =>  fabric_fpga_araddr_axi_s1_o(3)
       , fabric_fpga_araddr_axi_s1_o5                =>  fabric_fpga_araddr_axi_s1_o(4)
       , fabric_fpga_araddr_axi_s1_o6                =>  fabric_fpga_araddr_axi_s1_o(5)
       , fabric_fpga_araddr_axi_s1_o7                =>  fabric_fpga_araddr_axi_s1_o(6)
       , fabric_fpga_araddr_axi_s1_o8                =>  fabric_fpga_araddr_axi_s1_o(7)
       , fabric_fpga_araddr_axi_s1_o9                =>  fabric_fpga_araddr_axi_s1_o(8)
       , fabric_fpga_araddr_axi_s1_o10               =>  fabric_fpga_araddr_axi_s1_o(9)
       , fabric_fpga_araddr_axi_s1_o11               =>  fabric_fpga_araddr_axi_s1_o(10)
       , fabric_fpga_araddr_axi_s1_o12               =>  fabric_fpga_araddr_axi_s1_o(11)
       , fabric_fpga_araddr_axi_s1_o13               =>  fabric_fpga_araddr_axi_s1_o(12)
       , fabric_fpga_araddr_axi_s1_o14               =>  fabric_fpga_araddr_axi_s1_o(13)
       , fabric_fpga_araddr_axi_s1_o15               =>  fabric_fpga_araddr_axi_s1_o(14)
       , fabric_fpga_araddr_axi_s1_o16               =>  fabric_fpga_araddr_axi_s1_o(15)
       , fabric_fpga_araddr_axi_s1_o17               =>  fabric_fpga_araddr_axi_s1_o(16)
       , fabric_fpga_araddr_axi_s1_o18               =>  fabric_fpga_araddr_axi_s1_o(17)
       , fabric_fpga_araddr_axi_s1_o19               =>  fabric_fpga_araddr_axi_s1_o(18)
       , fabric_fpga_araddr_axi_s1_o20               =>  fabric_fpga_araddr_axi_s1_o(19)
       , fabric_fpga_araddr_axi_s1_o21               =>  fabric_fpga_araddr_axi_s1_o(20)
       , fabric_fpga_araddr_axi_s1_o22               =>  fabric_fpga_araddr_axi_s1_o(21)
       , fabric_fpga_araddr_axi_s1_o23               =>  fabric_fpga_araddr_axi_s1_o(22)
       , fabric_fpga_araddr_axi_s1_o24               =>  fabric_fpga_araddr_axi_s1_o(23)
       , fabric_fpga_araddr_axi_s1_o25               =>  fabric_fpga_araddr_axi_s1_o(24)
       , fabric_fpga_araddr_axi_s1_o26               =>  fabric_fpga_araddr_axi_s1_o(25)
       , fabric_fpga_araddr_axi_s1_o27               =>  fabric_fpga_araddr_axi_s1_o(26)
       , fabric_fpga_araddr_axi_s1_o28               =>  fabric_fpga_araddr_axi_s1_o(27)
       , fabric_fpga_araddr_axi_s1_o29               =>  fabric_fpga_araddr_axi_s1_o(28)
       , fabric_fpga_araddr_axi_s1_o30               =>  fabric_fpga_araddr_axi_s1_o(29)
       , fabric_fpga_araddr_axi_s1_o31               =>  fabric_fpga_araddr_axi_s1_o(30)
       , fabric_fpga_araddr_axi_s1_o32               =>  fabric_fpga_araddr_axi_s1_o(31)
       , fabric_fpga_araddr_axi_s1_o33               =>  fabric_fpga_araddr_axi_s1_o(32)
       , fabric_fpga_araddr_axi_s1_o34               =>  fabric_fpga_araddr_axi_s1_o(33)
       , fabric_fpga_araddr_axi_s1_o35               =>  fabric_fpga_araddr_axi_s1_o(34)
       , fabric_fpga_araddr_axi_s1_o36               =>  fabric_fpga_araddr_axi_s1_o(35)
       , fabric_fpga_araddr_axi_s1_o37               =>  fabric_fpga_araddr_axi_s1_o(36)
       , fabric_fpga_araddr_axi_s1_o38               =>  fabric_fpga_araddr_axi_s1_o(37)
       , fabric_fpga_araddr_axi_s1_o39               =>  fabric_fpga_araddr_axi_s1_o(38)
       , fabric_fpga_araddr_axi_s1_o40               =>  fabric_fpga_araddr_axi_s1_o(39)
       , fabric_fpga_arburst_axi_s1_o1               =>  fabric_fpga_arburst_axi_s1_o(0)
       , fabric_fpga_arburst_axi_s1_o2               =>  fabric_fpga_arburst_axi_s1_o(1)
       , fabric_fpga_arcache_axi_s1_o1               =>  fabric_fpga_arcache_axi_s1_o(0)
       , fabric_fpga_arcache_axi_s1_o2               =>  fabric_fpga_arcache_axi_s1_o(1)
       , fabric_fpga_arcache_axi_s1_o3               =>  fabric_fpga_arcache_axi_s1_o(2)
       , fabric_fpga_arcache_axi_s1_o4               =>  fabric_fpga_arcache_axi_s1_o(3)
       , fabric_fpga_arid_axi_s1_o1                  =>  fabric_fpga_arid_axi_s1_o(0)
       , fabric_fpga_arid_axi_s1_o2                  =>  fabric_fpga_arid_axi_s1_o(1)
       , fabric_fpga_arid_axi_s1_o3                  =>  fabric_fpga_arid_axi_s1_o(2)
       , fabric_fpga_arid_axi_s1_o4                  =>  fabric_fpga_arid_axi_s1_o(3)
       , fabric_fpga_arid_axi_s1_o5                  =>  fabric_fpga_arid_axi_s1_o(4)
       , fabric_fpga_arid_axi_s1_o6                  =>  fabric_fpga_arid_axi_s1_o(5)
       , fabric_fpga_arid_axi_s1_o7                  =>  fabric_fpga_arid_axi_s1_o(6)
       , fabric_fpga_arid_axi_s1_o8                  =>  fabric_fpga_arid_axi_s1_o(7)
       , fabric_fpga_arid_axi_s1_o9                  =>  fabric_fpga_arid_axi_s1_o(8)
       , fabric_fpga_arid_axi_s1_o10                 =>  fabric_fpga_arid_axi_s1_o(9)
       , fabric_fpga_arid_axi_s1_o11                 =>  fabric_fpga_arid_axi_s1_o(10)
       , fabric_fpga_arid_axi_s1_o12                 =>  fabric_fpga_arid_axi_s1_o(11)
       , fabric_fpga_arlen_axi_s1_o1                 =>  fabric_fpga_arlen_axi_s1_o(0)
       , fabric_fpga_arlen_axi_s1_o2                 =>  fabric_fpga_arlen_axi_s1_o(1)
       , fabric_fpga_arlen_axi_s1_o3                 =>  fabric_fpga_arlen_axi_s1_o(2)
       , fabric_fpga_arlen_axi_s1_o4                 =>  fabric_fpga_arlen_axi_s1_o(3)
       , fabric_fpga_arlen_axi_s1_o5                 =>  fabric_fpga_arlen_axi_s1_o(4)
       , fabric_fpga_arlen_axi_s1_o6                 =>  fabric_fpga_arlen_axi_s1_o(5)
       , fabric_fpga_arlen_axi_s1_o7                 =>  fabric_fpga_arlen_axi_s1_o(6)
       , fabric_fpga_arlen_axi_s1_o8                 =>  fabric_fpga_arlen_axi_s1_o(7)
       , fabric_fpga_arlock_axi_s1_o                 =>  fabric_fpga_arlock_axi_s1_o
       , fabric_fpga_arprot_axi_s1_o1                =>  fabric_fpga_arprot_axi_s1_o(0)
       , fabric_fpga_arprot_axi_s1_o2                =>  fabric_fpga_arprot_axi_s1_o(1)
       , fabric_fpga_arprot_axi_s1_o3                =>  fabric_fpga_arprot_axi_s1_o(2)
       , fabric_fpga_arqos_axi_s1_o1                 =>  fabric_fpga_arqos_axi_s1_o(0)
       , fabric_fpga_arqos_axi_s1_o2                 =>  fabric_fpga_arqos_axi_s1_o(1)
       , fabric_fpga_arqos_axi_s1_o3                 =>  fabric_fpga_arqos_axi_s1_o(2)
       , fabric_fpga_arqos_axi_s1_o4                 =>  fabric_fpga_arqos_axi_s1_o(3)
       , fabric_fpga_arregion_axi_s1_o1              =>  fabric_fpga_arregion_axi_s1_o(0)
       , fabric_fpga_arregion_axi_s1_o2              =>  fabric_fpga_arregion_axi_s1_o(1)
       , fabric_fpga_arregion_axi_s1_o3              =>  fabric_fpga_arregion_axi_s1_o(2)
       , fabric_fpga_arregion_axi_s1_o4              =>  fabric_fpga_arregion_axi_s1_o(3)
       , fabric_fpga_arsize_axi_s1_o1                =>  fabric_fpga_arsize_axi_s1_o(0)
       , fabric_fpga_arsize_axi_s1_o2                =>  fabric_fpga_arsize_axi_s1_o(1)
       , fabric_fpga_arsize_axi_s1_o3                =>  fabric_fpga_arsize_axi_s1_o(2)
       , fabric_fpga_arvalid_axi_s1_o                =>  fabric_fpga_arvalid_axi_s1_o
       , fabric_fpga_awaddr_axi_s1_o1                =>  fabric_fpga_awaddr_axi_s1_o(0)
       , fabric_fpga_awaddr_axi_s1_o2                =>  fabric_fpga_awaddr_axi_s1_o(1)
       , fabric_fpga_awaddr_axi_s1_o3                =>  fabric_fpga_awaddr_axi_s1_o(2)
       , fabric_fpga_awaddr_axi_s1_o4                =>  fabric_fpga_awaddr_axi_s1_o(3)
       , fabric_fpga_awaddr_axi_s1_o5                =>  fabric_fpga_awaddr_axi_s1_o(4)
       , fabric_fpga_awaddr_axi_s1_o6                =>  fabric_fpga_awaddr_axi_s1_o(5)
       , fabric_fpga_awaddr_axi_s1_o7                =>  fabric_fpga_awaddr_axi_s1_o(6)
       , fabric_fpga_awaddr_axi_s1_o8                =>  fabric_fpga_awaddr_axi_s1_o(7)
       , fabric_fpga_awaddr_axi_s1_o9                =>  fabric_fpga_awaddr_axi_s1_o(8)
       , fabric_fpga_awaddr_axi_s1_o10               =>  fabric_fpga_awaddr_axi_s1_o(9)
       , fabric_fpga_awaddr_axi_s1_o11               =>  fabric_fpga_awaddr_axi_s1_o(10)
       , fabric_fpga_awaddr_axi_s1_o12               =>  fabric_fpga_awaddr_axi_s1_o(11)
       , fabric_fpga_awaddr_axi_s1_o13               =>  fabric_fpga_awaddr_axi_s1_o(12)
       , fabric_fpga_awaddr_axi_s1_o14               =>  fabric_fpga_awaddr_axi_s1_o(13)
       , fabric_fpga_awaddr_axi_s1_o15               =>  fabric_fpga_awaddr_axi_s1_o(14)
       , fabric_fpga_awaddr_axi_s1_o16               =>  fabric_fpga_awaddr_axi_s1_o(15)
       , fabric_fpga_awaddr_axi_s1_o17               =>  fabric_fpga_awaddr_axi_s1_o(16)
       , fabric_fpga_awaddr_axi_s1_o18               =>  fabric_fpga_awaddr_axi_s1_o(17)
       , fabric_fpga_awaddr_axi_s1_o19               =>  fabric_fpga_awaddr_axi_s1_o(18)
       , fabric_fpga_awaddr_axi_s1_o20               =>  fabric_fpga_awaddr_axi_s1_o(19)
       , fabric_fpga_awaddr_axi_s1_o21               =>  fabric_fpga_awaddr_axi_s1_o(20)
       , fabric_fpga_awaddr_axi_s1_o22               =>  fabric_fpga_awaddr_axi_s1_o(21)
       , fabric_fpga_awaddr_axi_s1_o23               =>  fabric_fpga_awaddr_axi_s1_o(22)
       , fabric_fpga_awaddr_axi_s1_o24               =>  fabric_fpga_awaddr_axi_s1_o(23)
       , fabric_fpga_awaddr_axi_s1_o25               =>  fabric_fpga_awaddr_axi_s1_o(24)
       , fabric_fpga_awaddr_axi_s1_o26               =>  fabric_fpga_awaddr_axi_s1_o(25)
       , fabric_fpga_awaddr_axi_s1_o27               =>  fabric_fpga_awaddr_axi_s1_o(26)
       , fabric_fpga_awaddr_axi_s1_o28               =>  fabric_fpga_awaddr_axi_s1_o(27)
       , fabric_fpga_awaddr_axi_s1_o29               =>  fabric_fpga_awaddr_axi_s1_o(28)
       , fabric_fpga_awaddr_axi_s1_o30               =>  fabric_fpga_awaddr_axi_s1_o(29)
       , fabric_fpga_awaddr_axi_s1_o31               =>  fabric_fpga_awaddr_axi_s1_o(30)
       , fabric_fpga_awaddr_axi_s1_o32               =>  fabric_fpga_awaddr_axi_s1_o(31)
       , fabric_fpga_awaddr_axi_s1_o33               =>  fabric_fpga_awaddr_axi_s1_o(32)
       , fabric_fpga_awaddr_axi_s1_o34               =>  fabric_fpga_awaddr_axi_s1_o(33)
       , fabric_fpga_awaddr_axi_s1_o35               =>  fabric_fpga_awaddr_axi_s1_o(34)
       , fabric_fpga_awaddr_axi_s1_o36               =>  fabric_fpga_awaddr_axi_s1_o(35)
       , fabric_fpga_awaddr_axi_s1_o37               =>  fabric_fpga_awaddr_axi_s1_o(36)
       , fabric_fpga_awaddr_axi_s1_o38               =>  fabric_fpga_awaddr_axi_s1_o(37)
       , fabric_fpga_awaddr_axi_s1_o39               =>  fabric_fpga_awaddr_axi_s1_o(38)
       , fabric_fpga_awaddr_axi_s1_o40               =>  fabric_fpga_awaddr_axi_s1_o(39)
       , fabric_fpga_awburst_axi_s1_o1               =>  fabric_fpga_awburst_axi_s1_o(0)
       , fabric_fpga_awburst_axi_s1_o2               =>  fabric_fpga_awburst_axi_s1_o(1)
       , fabric_fpga_awcache_axi_s1_o1               =>  fabric_fpga_awcache_axi_s1_o(0)
       , fabric_fpga_awcache_axi_s1_o2               =>  fabric_fpga_awcache_axi_s1_o(1)
       , fabric_fpga_awcache_axi_s1_o3               =>  fabric_fpga_awcache_axi_s1_o(2)
       , fabric_fpga_awcache_axi_s1_o4               =>  fabric_fpga_awcache_axi_s1_o(3)
       , fabric_fpga_awid_axi_s1_o1                  =>  fabric_fpga_awid_axi_s1_o(0)
       , fabric_fpga_awid_axi_s1_o2                  =>  fabric_fpga_awid_axi_s1_o(1)
       , fabric_fpga_awid_axi_s1_o3                  =>  fabric_fpga_awid_axi_s1_o(2)
       , fabric_fpga_awid_axi_s1_o4                  =>  fabric_fpga_awid_axi_s1_o(3)
       , fabric_fpga_awid_axi_s1_o5                  =>  fabric_fpga_awid_axi_s1_o(4)
       , fabric_fpga_awid_axi_s1_o6                  =>  fabric_fpga_awid_axi_s1_o(5)
       , fabric_fpga_awid_axi_s1_o7                  =>  fabric_fpga_awid_axi_s1_o(6)
       , fabric_fpga_awid_axi_s1_o8                  =>  fabric_fpga_awid_axi_s1_o(7)
       , fabric_fpga_awid_axi_s1_o9                  =>  fabric_fpga_awid_axi_s1_o(8)
       , fabric_fpga_awid_axi_s1_o10                 =>  fabric_fpga_awid_axi_s1_o(9)
       , fabric_fpga_awid_axi_s1_o11                 =>  fabric_fpga_awid_axi_s1_o(10)
       , fabric_fpga_awid_axi_s1_o12                 =>  fabric_fpga_awid_axi_s1_o(11)
       , fabric_fpga_awlen_axi_s1_o1                 =>  fabric_fpga_awlen_axi_s1_o(0)
       , fabric_fpga_awlen_axi_s1_o2                 =>  fabric_fpga_awlen_axi_s1_o(1)
       , fabric_fpga_awlen_axi_s1_o3                 =>  fabric_fpga_awlen_axi_s1_o(2)
       , fabric_fpga_awlen_axi_s1_o4                 =>  fabric_fpga_awlen_axi_s1_o(3)
       , fabric_fpga_awlen_axi_s1_o5                 =>  fabric_fpga_awlen_axi_s1_o(4)
       , fabric_fpga_awlen_axi_s1_o6                 =>  fabric_fpga_awlen_axi_s1_o(5)
       , fabric_fpga_awlen_axi_s1_o7                 =>  fabric_fpga_awlen_axi_s1_o(6)
       , fabric_fpga_awlen_axi_s1_o8                 =>  fabric_fpga_awlen_axi_s1_o(7)
       , fabric_fpga_awlock_axi_s1_o                 =>  fabric_fpga_awlock_axi_s1_o
       , fabric_fpga_awprot_axi_s1_o1                =>  fabric_fpga_awprot_axi_s1_o(0)
       , fabric_fpga_awprot_axi_s1_o2                =>  fabric_fpga_awprot_axi_s1_o(1)
       , fabric_fpga_awprot_axi_s1_o3                =>  fabric_fpga_awprot_axi_s1_o(2)
       , fabric_fpga_awqos_axi_s1_o1                 =>  fabric_fpga_awqos_axi_s1_o(0)
       , fabric_fpga_awqos_axi_s1_o2                 =>  fabric_fpga_awqos_axi_s1_o(1)
       , fabric_fpga_awqos_axi_s1_o3                 =>  fabric_fpga_awqos_axi_s1_o(2)
       , fabric_fpga_awqos_axi_s1_o4                 =>  fabric_fpga_awqos_axi_s1_o(3)
       , fabric_fpga_awregion_axi_s1_o1              =>  fabric_fpga_awregion_axi_s1_o(0)
       , fabric_fpga_awregion_axi_s1_o2              =>  fabric_fpga_awregion_axi_s1_o(1)
       , fabric_fpga_awregion_axi_s1_o3              =>  fabric_fpga_awregion_axi_s1_o(2)
       , fabric_fpga_awregion_axi_s1_o4              =>  fabric_fpga_awregion_axi_s1_o(3)
       , fabric_fpga_awsize_axi_s1_o1                =>  fabric_fpga_awsize_axi_s1_o(0)
       , fabric_fpga_awsize_axi_s1_o2                =>  fabric_fpga_awsize_axi_s1_o(1)
       , fabric_fpga_awsize_axi_s1_o3                =>  fabric_fpga_awsize_axi_s1_o(2)
       , fabric_fpga_bready_axi_s1_o                 =>  fabric_fpga_bready_axi_s1_o
       , fabric_fpga_rready_axi_s1_o                 =>  fabric_fpga_rready_axi_s1_o
       , fabric_fpga_wdata_axi_s1_o1                 =>  fabric_fpga_wdata_axi_s1_o(0)
       , fabric_fpga_wdata_axi_s1_o2                 =>  fabric_fpga_wdata_axi_s1_o(1)
       , fabric_fpga_wdata_axi_s1_o3                 =>  fabric_fpga_wdata_axi_s1_o(2)
       , fabric_fpga_wdata_axi_s1_o4                 =>  fabric_fpga_wdata_axi_s1_o(3)
       , fabric_fpga_wdata_axi_s1_o5                 =>  fabric_fpga_wdata_axi_s1_o(4)
       , fabric_fpga_wdata_axi_s1_o6                 =>  fabric_fpga_wdata_axi_s1_o(5)
       , fabric_fpga_wdata_axi_s1_o7                 =>  fabric_fpga_wdata_axi_s1_o(6)
       , fabric_fpga_wdata_axi_s1_o8                 =>  fabric_fpga_wdata_axi_s1_o(7)
       , fabric_fpga_wdata_axi_s1_o9                 =>  fabric_fpga_wdata_axi_s1_o(8)
       , fabric_fpga_wdata_axi_s1_o10                =>  fabric_fpga_wdata_axi_s1_o(9)
       , fabric_fpga_wdata_axi_s1_o11                =>  fabric_fpga_wdata_axi_s1_o(10)
       , fabric_fpga_wdata_axi_s1_o12                =>  fabric_fpga_wdata_axi_s1_o(11)
       , fabric_fpga_wdata_axi_s1_o13                =>  fabric_fpga_wdata_axi_s1_o(12)
       , fabric_fpga_wdata_axi_s1_o14                =>  fabric_fpga_wdata_axi_s1_o(13)
       , fabric_fpga_wdata_axi_s1_o15                =>  fabric_fpga_wdata_axi_s1_o(14)
       , fabric_fpga_wdata_axi_s1_o16                =>  fabric_fpga_wdata_axi_s1_o(15)
       , fabric_fpga_wdata_axi_s1_o17                =>  fabric_fpga_wdata_axi_s1_o(16)
       , fabric_fpga_wdata_axi_s1_o18                =>  fabric_fpga_wdata_axi_s1_o(17)
       , fabric_fpga_wdata_axi_s1_o19                =>  fabric_fpga_wdata_axi_s1_o(18)
       , fabric_fpga_wdata_axi_s1_o20                =>  fabric_fpga_wdata_axi_s1_o(19)
       , fabric_fpga_wdata_axi_s1_o21                =>  fabric_fpga_wdata_axi_s1_o(20)
       , fabric_fpga_wdata_axi_s1_o22                =>  fabric_fpga_wdata_axi_s1_o(21)
       , fabric_fpga_wdata_axi_s1_o23                =>  fabric_fpga_wdata_axi_s1_o(22)
       , fabric_fpga_wdata_axi_s1_o24                =>  fabric_fpga_wdata_axi_s1_o(23)
       , fabric_fpga_wdata_axi_s1_o25                =>  fabric_fpga_wdata_axi_s1_o(24)
       , fabric_fpga_wdata_axi_s1_o26                =>  fabric_fpga_wdata_axi_s1_o(25)
       , fabric_fpga_wdata_axi_s1_o27                =>  fabric_fpga_wdata_axi_s1_o(26)
       , fabric_fpga_wdata_axi_s1_o28                =>  fabric_fpga_wdata_axi_s1_o(27)
       , fabric_fpga_wdata_axi_s1_o29                =>  fabric_fpga_wdata_axi_s1_o(28)
       , fabric_fpga_wdata_axi_s1_o30                =>  fabric_fpga_wdata_axi_s1_o(29)
       , fabric_fpga_wdata_axi_s1_o31                =>  fabric_fpga_wdata_axi_s1_o(30)
       , fabric_fpga_wdata_axi_s1_o32                =>  fabric_fpga_wdata_axi_s1_o(31)
       , fabric_fpga_wdata_axi_s1_o33                =>  fabric_fpga_wdata_axi_s1_o(32)
       , fabric_fpga_wdata_axi_s1_o34                =>  fabric_fpga_wdata_axi_s1_o(33)
       , fabric_fpga_wdata_axi_s1_o35                =>  fabric_fpga_wdata_axi_s1_o(34)
       , fabric_fpga_wdata_axi_s1_o36                =>  fabric_fpga_wdata_axi_s1_o(35)
       , fabric_fpga_wdata_axi_s1_o37                =>  fabric_fpga_wdata_axi_s1_o(36)
       , fabric_fpga_wdata_axi_s1_o38                =>  fabric_fpga_wdata_axi_s1_o(37)
       , fabric_fpga_wdata_axi_s1_o39                =>  fabric_fpga_wdata_axi_s1_o(38)
       , fabric_fpga_wdata_axi_s1_o40                =>  fabric_fpga_wdata_axi_s1_o(39)
       , fabric_fpga_wdata_axi_s1_o41                =>  fabric_fpga_wdata_axi_s1_o(40)
       , fabric_fpga_wdata_axi_s1_o42                =>  fabric_fpga_wdata_axi_s1_o(41)
       , fabric_fpga_wdata_axi_s1_o43                =>  fabric_fpga_wdata_axi_s1_o(42)
       , fabric_fpga_wdata_axi_s1_o44                =>  fabric_fpga_wdata_axi_s1_o(43)
       , fabric_fpga_wdata_axi_s1_o45                =>  fabric_fpga_wdata_axi_s1_o(44)
       , fabric_fpga_wdata_axi_s1_o46                =>  fabric_fpga_wdata_axi_s1_o(45)
       , fabric_fpga_wdata_axi_s1_o47                =>  fabric_fpga_wdata_axi_s1_o(46)
       , fabric_fpga_wdata_axi_s1_o48                =>  fabric_fpga_wdata_axi_s1_o(47)
       , fabric_fpga_wdata_axi_s1_o49                =>  fabric_fpga_wdata_axi_s1_o(48)
       , fabric_fpga_wdata_axi_s1_o50                =>  fabric_fpga_wdata_axi_s1_o(49)
       , fabric_fpga_wdata_axi_s1_o51                =>  fabric_fpga_wdata_axi_s1_o(50)
       , fabric_fpga_wdata_axi_s1_o52                =>  fabric_fpga_wdata_axi_s1_o(51)
       , fabric_fpga_wdata_axi_s1_o53                =>  fabric_fpga_wdata_axi_s1_o(52)
       , fabric_fpga_wdata_axi_s1_o54                =>  fabric_fpga_wdata_axi_s1_o(53)
       , fabric_fpga_wdata_axi_s1_o55                =>  fabric_fpga_wdata_axi_s1_o(54)
       , fabric_fpga_wdata_axi_s1_o56                =>  fabric_fpga_wdata_axi_s1_o(55)
       , fabric_fpga_wdata_axi_s1_o57                =>  fabric_fpga_wdata_axi_s1_o(56)
       , fabric_fpga_wdata_axi_s1_o58                =>  fabric_fpga_wdata_axi_s1_o(57)
       , fabric_fpga_wdata_axi_s1_o59                =>  fabric_fpga_wdata_axi_s1_o(58)
       , fabric_fpga_wdata_axi_s1_o60                =>  fabric_fpga_wdata_axi_s1_o(59)
       , fabric_fpga_wdata_axi_s1_o61                =>  fabric_fpga_wdata_axi_s1_o(60)
       , fabric_fpga_wdata_axi_s1_o62                =>  fabric_fpga_wdata_axi_s1_o(61)
       , fabric_fpga_wdata_axi_s1_o63                =>  fabric_fpga_wdata_axi_s1_o(62)
       , fabric_fpga_wdata_axi_s1_o64                =>  fabric_fpga_wdata_axi_s1_o(63)
       , fabric_fpga_wdata_axi_s1_o65                =>  fabric_fpga_wdata_axi_s1_o(64)
       , fabric_fpga_wdata_axi_s1_o66                =>  fabric_fpga_wdata_axi_s1_o(65)
       , fabric_fpga_wdata_axi_s1_o67                =>  fabric_fpga_wdata_axi_s1_o(66)
       , fabric_fpga_wdata_axi_s1_o68                =>  fabric_fpga_wdata_axi_s1_o(67)
       , fabric_fpga_wdata_axi_s1_o69                =>  fabric_fpga_wdata_axi_s1_o(68)
       , fabric_fpga_wdata_axi_s1_o70                =>  fabric_fpga_wdata_axi_s1_o(69)
       , fabric_fpga_wdata_axi_s1_o71                =>  fabric_fpga_wdata_axi_s1_o(70)
       , fabric_fpga_wdata_axi_s1_o72                =>  fabric_fpga_wdata_axi_s1_o(71)
       , fabric_fpga_wdata_axi_s1_o73                =>  fabric_fpga_wdata_axi_s1_o(72)
       , fabric_fpga_wdata_axi_s1_o74                =>  fabric_fpga_wdata_axi_s1_o(73)
       , fabric_fpga_wdata_axi_s1_o75                =>  fabric_fpga_wdata_axi_s1_o(74)
       , fabric_fpga_wdata_axi_s1_o76                =>  fabric_fpga_wdata_axi_s1_o(75)
       , fabric_fpga_wdata_axi_s1_o77                =>  fabric_fpga_wdata_axi_s1_o(76)
       , fabric_fpga_wdata_axi_s1_o78                =>  fabric_fpga_wdata_axi_s1_o(77)
       , fabric_fpga_wdata_axi_s1_o79                =>  fabric_fpga_wdata_axi_s1_o(78)
       , fabric_fpga_wdata_axi_s1_o80                =>  fabric_fpga_wdata_axi_s1_o(79)
       , fabric_fpga_wdata_axi_s1_o81                =>  fabric_fpga_wdata_axi_s1_o(80)
       , fabric_fpga_wdata_axi_s1_o82                =>  fabric_fpga_wdata_axi_s1_o(81)
       , fabric_fpga_wdata_axi_s1_o83                =>  fabric_fpga_wdata_axi_s1_o(82)
       , fabric_fpga_wdata_axi_s1_o84                =>  fabric_fpga_wdata_axi_s1_o(83)
       , fabric_fpga_wdata_axi_s1_o85                =>  fabric_fpga_wdata_axi_s1_o(84)
       , fabric_fpga_wdata_axi_s1_o86                =>  fabric_fpga_wdata_axi_s1_o(85)
       , fabric_fpga_wdata_axi_s1_o87                =>  fabric_fpga_wdata_axi_s1_o(86)
       , fabric_fpga_wdata_axi_s1_o88                =>  fabric_fpga_wdata_axi_s1_o(87)
       , fabric_fpga_wdata_axi_s1_o89                =>  fabric_fpga_wdata_axi_s1_o(88)
       , fabric_fpga_wdata_axi_s1_o90                =>  fabric_fpga_wdata_axi_s1_o(89)
       , fabric_fpga_wdata_axi_s1_o91                =>  fabric_fpga_wdata_axi_s1_o(90)
       , fabric_fpga_wdata_axi_s1_o92                =>  fabric_fpga_wdata_axi_s1_o(91)
       , fabric_fpga_wdata_axi_s1_o93                =>  fabric_fpga_wdata_axi_s1_o(92)
       , fabric_fpga_wdata_axi_s1_o94                =>  fabric_fpga_wdata_axi_s1_o(93)
       , fabric_fpga_wdata_axi_s1_o95                =>  fabric_fpga_wdata_axi_s1_o(94)
       , fabric_fpga_wdata_axi_s1_o96                =>  fabric_fpga_wdata_axi_s1_o(95)
       , fabric_fpga_wdata_axi_s1_o97                =>  fabric_fpga_wdata_axi_s1_o(96)
       , fabric_fpga_wdata_axi_s1_o98                =>  fabric_fpga_wdata_axi_s1_o(97)
       , fabric_fpga_wdata_axi_s1_o99                =>  fabric_fpga_wdata_axi_s1_o(98)
       , fabric_fpga_wdata_axi_s1_o100               =>  fabric_fpga_wdata_axi_s1_o(99)
       , fabric_fpga_wdata_axi_s1_o101               =>  fabric_fpga_wdata_axi_s1_o(100)
       , fabric_fpga_wdata_axi_s1_o102               =>  fabric_fpga_wdata_axi_s1_o(101)
       , fabric_fpga_wdata_axi_s1_o103               =>  fabric_fpga_wdata_axi_s1_o(102)
       , fabric_fpga_wdata_axi_s1_o104               =>  fabric_fpga_wdata_axi_s1_o(103)
       , fabric_fpga_wdata_axi_s1_o105               =>  fabric_fpga_wdata_axi_s1_o(104)
       , fabric_fpga_wdata_axi_s1_o106               =>  fabric_fpga_wdata_axi_s1_o(105)
       , fabric_fpga_wdata_axi_s1_o107               =>  fabric_fpga_wdata_axi_s1_o(106)
       , fabric_fpga_wdata_axi_s1_o108               =>  fabric_fpga_wdata_axi_s1_o(107)
       , fabric_fpga_wdata_axi_s1_o109               =>  fabric_fpga_wdata_axi_s1_o(108)
       , fabric_fpga_wdata_axi_s1_o110               =>  fabric_fpga_wdata_axi_s1_o(109)
       , fabric_fpga_wdata_axi_s1_o111               =>  fabric_fpga_wdata_axi_s1_o(110)
       , fabric_fpga_wdata_axi_s1_o112               =>  fabric_fpga_wdata_axi_s1_o(111)
       , fabric_fpga_wdata_axi_s1_o113               =>  fabric_fpga_wdata_axi_s1_o(112)
       , fabric_fpga_wdata_axi_s1_o114               =>  fabric_fpga_wdata_axi_s1_o(113)
       , fabric_fpga_wdata_axi_s1_o115               =>  fabric_fpga_wdata_axi_s1_o(114)
       , fabric_fpga_wdata_axi_s1_o116               =>  fabric_fpga_wdata_axi_s1_o(115)
       , fabric_fpga_wdata_axi_s1_o117               =>  fabric_fpga_wdata_axi_s1_o(116)
       , fabric_fpga_wdata_axi_s1_o118               =>  fabric_fpga_wdata_axi_s1_o(117)
       , fabric_fpga_wdata_axi_s1_o119               =>  fabric_fpga_wdata_axi_s1_o(118)
       , fabric_fpga_wdata_axi_s1_o120               =>  fabric_fpga_wdata_axi_s1_o(119)
       , fabric_fpga_wdata_axi_s1_o121               =>  fabric_fpga_wdata_axi_s1_o(120)
       , fabric_fpga_wdata_axi_s1_o122               =>  fabric_fpga_wdata_axi_s1_o(121)
       , fabric_fpga_wdata_axi_s1_o123               =>  fabric_fpga_wdata_axi_s1_o(122)
       , fabric_fpga_wdata_axi_s1_o124               =>  fabric_fpga_wdata_axi_s1_o(123)
       , fabric_fpga_wdata_axi_s1_o125               =>  fabric_fpga_wdata_axi_s1_o(124)
       , fabric_fpga_wdata_axi_s1_o126               =>  fabric_fpga_wdata_axi_s1_o(125)
       , fabric_fpga_wdata_axi_s1_o127               =>  fabric_fpga_wdata_axi_s1_o(126)
       , fabric_fpga_wdata_axi_s1_o128               =>  fabric_fpga_wdata_axi_s1_o(127)
       , fabric_fpga_wlast_axi_s1_o                  =>  fabric_fpga_wlast_axi_s1_o
       , fabric_fpga_wstrb_axi_s1_o1                 =>  fabric_fpga_wstrb_axi_s1_o(0)
       , fabric_fpga_wstrb_axi_s1_o2                 =>  fabric_fpga_wstrb_axi_s1_o(1)
       , fabric_fpga_wstrb_axi_s1_o3                 =>  fabric_fpga_wstrb_axi_s1_o(2)
       , fabric_fpga_wstrb_axi_s1_o4                 =>  fabric_fpga_wstrb_axi_s1_o(3)
       , fabric_fpga_wstrb_axi_s1_o5                 =>  fabric_fpga_wstrb_axi_s1_o(4)
       , fabric_fpga_wstrb_axi_s1_o6                 =>  fabric_fpga_wstrb_axi_s1_o(5)
       , fabric_fpga_wstrb_axi_s1_o7                 =>  fabric_fpga_wstrb_axi_s1_o(6)
       , fabric_fpga_wstrb_axi_s1_o8                 =>  fabric_fpga_wstrb_axi_s1_o(7)
       , fabric_fpga_wstrb_axi_s1_o9                 =>  fabric_fpga_wstrb_axi_s1_o(8)
       , fabric_fpga_wstrb_axi_s1_o10                =>  fabric_fpga_wstrb_axi_s1_o(9)
       , fabric_fpga_wstrb_axi_s1_o11                =>  fabric_fpga_wstrb_axi_s1_o(10)
       , fabric_fpga_wstrb_axi_s1_o12                =>  fabric_fpga_wstrb_axi_s1_o(11)
       , fabric_fpga_wstrb_axi_s1_o13                =>  fabric_fpga_wstrb_axi_s1_o(12)
       , fabric_fpga_wstrb_axi_s1_o14                =>  fabric_fpga_wstrb_axi_s1_o(13)
       , fabric_fpga_wstrb_axi_s1_o15                =>  fabric_fpga_wstrb_axi_s1_o(14)
       , fabric_fpga_wstrb_axi_s1_o16                =>  fabric_fpga_wstrb_axi_s1_o(15)
       , fabric_fpga_wvalid_axi_s1_o                 =>  fabric_fpga_wvalid_axi_s1_o
       , fabric_fpga_awvalid_axi_s1_o                =>  fabric_fpga_awvalid_axi_s1_o
       , fabric_fpga_arready_axi_s1_i                =>  fabric_fpga_arready_axi_s1_i
       , fabric_fpga_awready_axi_s1_i                =>  fabric_fpga_awready_axi_s1_i
       , fabric_fpga_bid_axi_s1_i1                   =>  fabric_fpga_bid_axi_s1_i(0)
       , fabric_fpga_bid_axi_s1_i2                   =>  fabric_fpga_bid_axi_s1_i(1)
       , fabric_fpga_bid_axi_s1_i3                   =>  fabric_fpga_bid_axi_s1_i(2)
       , fabric_fpga_bid_axi_s1_i4                   =>  fabric_fpga_bid_axi_s1_i(3)
       , fabric_fpga_bid_axi_s1_i5                   =>  fabric_fpga_bid_axi_s1_i(4)
       , fabric_fpga_bid_axi_s1_i6                   =>  fabric_fpga_bid_axi_s1_i(5)
       , fabric_fpga_bid_axi_s1_i7                   =>  fabric_fpga_bid_axi_s1_i(6)
       , fabric_fpga_bid_axi_s1_i8                   =>  fabric_fpga_bid_axi_s1_i(7)
       , fabric_fpga_bid_axi_s1_i9                   =>  fabric_fpga_bid_axi_s1_i(8)
       , fabric_fpga_bid_axi_s1_i10                  =>  fabric_fpga_bid_axi_s1_i(9)
       , fabric_fpga_bid_axi_s1_i11                  =>  fabric_fpga_bid_axi_s1_i(10)
       , fabric_fpga_bid_axi_s1_i12                  =>  fabric_fpga_bid_axi_s1_i(11)
       , fabric_fpga_bresp_axi_s1_i1                 =>  fabric_fpga_bresp_axi_s1_i(0)
       , fabric_fpga_bresp_axi_s1_i2                 =>  fabric_fpga_bresp_axi_s1_i(1)
       , fabric_fpga_bvalid_axi_s1_i                 =>  fabric_fpga_bvalid_axi_s1_i
       , fabric_fpga_rdata_axi_s1_i1                 =>  fabric_fpga_rdata_axi_s1_i(0)
       , fabric_fpga_rdata_axi_s1_i2                 =>  fabric_fpga_rdata_axi_s1_i(1)
       , fabric_fpga_rdata_axi_s1_i3                 =>  fabric_fpga_rdata_axi_s1_i(2)
       , fabric_fpga_rdata_axi_s1_i4                 =>  fabric_fpga_rdata_axi_s1_i(3)
       , fabric_fpga_rdata_axi_s1_i5                 =>  fabric_fpga_rdata_axi_s1_i(4)
       , fabric_fpga_rdata_axi_s1_i6                 =>  fabric_fpga_rdata_axi_s1_i(5)
       , fabric_fpga_rdata_axi_s1_i7                 =>  fabric_fpga_rdata_axi_s1_i(6)
       , fabric_fpga_rdata_axi_s1_i8                 =>  fabric_fpga_rdata_axi_s1_i(7)
       , fabric_fpga_rdata_axi_s1_i9                 =>  fabric_fpga_rdata_axi_s1_i(8)
       , fabric_fpga_rdata_axi_s1_i10                =>  fabric_fpga_rdata_axi_s1_i(9)
       , fabric_fpga_rdata_axi_s1_i11                =>  fabric_fpga_rdata_axi_s1_i(10)
       , fabric_fpga_rdata_axi_s1_i12                =>  fabric_fpga_rdata_axi_s1_i(11)
       , fabric_fpga_rdata_axi_s1_i13                =>  fabric_fpga_rdata_axi_s1_i(12)
       , fabric_fpga_rdata_axi_s1_i14                =>  fabric_fpga_rdata_axi_s1_i(13)
       , fabric_fpga_rdata_axi_s1_i15                =>  fabric_fpga_rdata_axi_s1_i(14)
       , fabric_fpga_rdata_axi_s1_i16                =>  fabric_fpga_rdata_axi_s1_i(15)
       , fabric_fpga_rdata_axi_s1_i17                =>  fabric_fpga_rdata_axi_s1_i(16)
       , fabric_fpga_rdata_axi_s1_i18                =>  fabric_fpga_rdata_axi_s1_i(17)
       , fabric_fpga_rdata_axi_s1_i19                =>  fabric_fpga_rdata_axi_s1_i(18)
       , fabric_fpga_rdata_axi_s1_i20                =>  fabric_fpga_rdata_axi_s1_i(19)
       , fabric_fpga_rdata_axi_s1_i21                =>  fabric_fpga_rdata_axi_s1_i(20)
       , fabric_fpga_rdata_axi_s1_i22                =>  fabric_fpga_rdata_axi_s1_i(21)
       , fabric_fpga_rdata_axi_s1_i23                =>  fabric_fpga_rdata_axi_s1_i(22)
       , fabric_fpga_rdata_axi_s1_i24                =>  fabric_fpga_rdata_axi_s1_i(23)
       , fabric_fpga_rdata_axi_s1_i25                =>  fabric_fpga_rdata_axi_s1_i(24)
       , fabric_fpga_rdata_axi_s1_i26                =>  fabric_fpga_rdata_axi_s1_i(25)
       , fabric_fpga_rdata_axi_s1_i27                =>  fabric_fpga_rdata_axi_s1_i(26)
       , fabric_fpga_rdata_axi_s1_i28                =>  fabric_fpga_rdata_axi_s1_i(27)
       , fabric_fpga_rdata_axi_s1_i29                =>  fabric_fpga_rdata_axi_s1_i(28)
       , fabric_fpga_rdata_axi_s1_i30                =>  fabric_fpga_rdata_axi_s1_i(29)
       , fabric_fpga_rdata_axi_s1_i31                =>  fabric_fpga_rdata_axi_s1_i(30)
       , fabric_fpga_rdata_axi_s1_i32                =>  fabric_fpga_rdata_axi_s1_i(31)
       , fabric_fpga_rdata_axi_s1_i33                =>  fabric_fpga_rdata_axi_s1_i(32)
       , fabric_fpga_rdata_axi_s1_i34                =>  fabric_fpga_rdata_axi_s1_i(33)
       , fabric_fpga_rdata_axi_s1_i35                =>  fabric_fpga_rdata_axi_s1_i(34)
       , fabric_fpga_rdata_axi_s1_i36                =>  fabric_fpga_rdata_axi_s1_i(35)
       , fabric_fpga_rdata_axi_s1_i37                =>  fabric_fpga_rdata_axi_s1_i(36)
       , fabric_fpga_rdata_axi_s1_i38                =>  fabric_fpga_rdata_axi_s1_i(37)
       , fabric_fpga_rdata_axi_s1_i39                =>  fabric_fpga_rdata_axi_s1_i(38)
       , fabric_fpga_rdata_axi_s1_i40                =>  fabric_fpga_rdata_axi_s1_i(39)
       , fabric_fpga_rdata_axi_s1_i41                =>  fabric_fpga_rdata_axi_s1_i(40)
       , fabric_fpga_rdata_axi_s1_i42                =>  fabric_fpga_rdata_axi_s1_i(41)
       , fabric_fpga_rdata_axi_s1_i43                =>  fabric_fpga_rdata_axi_s1_i(42)
       , fabric_fpga_rdata_axi_s1_i44                =>  fabric_fpga_rdata_axi_s1_i(43)
       , fabric_fpga_rdata_axi_s1_i45                =>  fabric_fpga_rdata_axi_s1_i(44)
       , fabric_fpga_rdata_axi_s1_i46                =>  fabric_fpga_rdata_axi_s1_i(45)
       , fabric_fpga_rdata_axi_s1_i47                =>  fabric_fpga_rdata_axi_s1_i(46)
       , fabric_fpga_rdata_axi_s1_i48                =>  fabric_fpga_rdata_axi_s1_i(47)
       , fabric_fpga_rdata_axi_s1_i49                =>  fabric_fpga_rdata_axi_s1_i(48)
       , fabric_fpga_rdata_axi_s1_i50                =>  fabric_fpga_rdata_axi_s1_i(49)
       , fabric_fpga_rdata_axi_s1_i51                =>  fabric_fpga_rdata_axi_s1_i(50)
       , fabric_fpga_rdata_axi_s1_i52                =>  fabric_fpga_rdata_axi_s1_i(51)
       , fabric_fpga_rdata_axi_s1_i53                =>  fabric_fpga_rdata_axi_s1_i(52)
       , fabric_fpga_rdata_axi_s1_i54                =>  fabric_fpga_rdata_axi_s1_i(53)
       , fabric_fpga_rdata_axi_s1_i55                =>  fabric_fpga_rdata_axi_s1_i(54)
       , fabric_fpga_rdata_axi_s1_i56                =>  fabric_fpga_rdata_axi_s1_i(55)
       , fabric_fpga_rdata_axi_s1_i57                =>  fabric_fpga_rdata_axi_s1_i(56)
       , fabric_fpga_rdata_axi_s1_i58                =>  fabric_fpga_rdata_axi_s1_i(57)
       , fabric_fpga_rdata_axi_s1_i59                =>  fabric_fpga_rdata_axi_s1_i(58)
       , fabric_fpga_rdata_axi_s1_i60                =>  fabric_fpga_rdata_axi_s1_i(59)
       , fabric_fpga_rdata_axi_s1_i61                =>  fabric_fpga_rdata_axi_s1_i(60)
       , fabric_fpga_rdata_axi_s1_i62                =>  fabric_fpga_rdata_axi_s1_i(61)
       , fabric_fpga_rdata_axi_s1_i63                =>  fabric_fpga_rdata_axi_s1_i(62)
       , fabric_fpga_rdata_axi_s1_i64                =>  fabric_fpga_rdata_axi_s1_i(63)
       , fabric_fpga_rdata_axi_s1_i65                =>  fabric_fpga_rdata_axi_s1_i(64)
       , fabric_fpga_rdata_axi_s1_i66                =>  fabric_fpga_rdata_axi_s1_i(65)
       , fabric_fpga_rdata_axi_s1_i67                =>  fabric_fpga_rdata_axi_s1_i(66)
       , fabric_fpga_rdata_axi_s1_i68                =>  fabric_fpga_rdata_axi_s1_i(67)
       , fabric_fpga_rdata_axi_s1_i69                =>  fabric_fpga_rdata_axi_s1_i(68)
       , fabric_fpga_rdata_axi_s1_i70                =>  fabric_fpga_rdata_axi_s1_i(69)
       , fabric_fpga_rdata_axi_s1_i71                =>  fabric_fpga_rdata_axi_s1_i(70)
       , fabric_fpga_rdata_axi_s1_i72                =>  fabric_fpga_rdata_axi_s1_i(71)
       , fabric_fpga_rdata_axi_s1_i73                =>  fabric_fpga_rdata_axi_s1_i(72)
       , fabric_fpga_rdata_axi_s1_i74                =>  fabric_fpga_rdata_axi_s1_i(73)
       , fabric_fpga_rdata_axi_s1_i75                =>  fabric_fpga_rdata_axi_s1_i(74)
       , fabric_fpga_rdata_axi_s1_i76                =>  fabric_fpga_rdata_axi_s1_i(75)
       , fabric_fpga_rdata_axi_s1_i77                =>  fabric_fpga_rdata_axi_s1_i(76)
       , fabric_fpga_rdata_axi_s1_i78                =>  fabric_fpga_rdata_axi_s1_i(77)
       , fabric_fpga_rdata_axi_s1_i79                =>  fabric_fpga_rdata_axi_s1_i(78)
       , fabric_fpga_rdata_axi_s1_i80                =>  fabric_fpga_rdata_axi_s1_i(79)
       , fabric_fpga_rdata_axi_s1_i81                =>  fabric_fpga_rdata_axi_s1_i(80)
       , fabric_fpga_rdata_axi_s1_i82                =>  fabric_fpga_rdata_axi_s1_i(81)
       , fabric_fpga_rdata_axi_s1_i83                =>  fabric_fpga_rdata_axi_s1_i(82)
       , fabric_fpga_rdata_axi_s1_i84                =>  fabric_fpga_rdata_axi_s1_i(83)
       , fabric_fpga_rdata_axi_s1_i85                =>  fabric_fpga_rdata_axi_s1_i(84)
       , fabric_fpga_rdata_axi_s1_i86                =>  fabric_fpga_rdata_axi_s1_i(85)
       , fabric_fpga_rdata_axi_s1_i87                =>  fabric_fpga_rdata_axi_s1_i(86)
       , fabric_fpga_rdata_axi_s1_i88                =>  fabric_fpga_rdata_axi_s1_i(87)
       , fabric_fpga_rdata_axi_s1_i89                =>  fabric_fpga_rdata_axi_s1_i(88)
       , fabric_fpga_rdata_axi_s1_i90                =>  fabric_fpga_rdata_axi_s1_i(89)
       , fabric_fpga_rdata_axi_s1_i91                =>  fabric_fpga_rdata_axi_s1_i(90)
       , fabric_fpga_rdata_axi_s1_i92                =>  fabric_fpga_rdata_axi_s1_i(91)
       , fabric_fpga_rdata_axi_s1_i93                =>  fabric_fpga_rdata_axi_s1_i(92)
       , fabric_fpga_rdata_axi_s1_i94                =>  fabric_fpga_rdata_axi_s1_i(93)
       , fabric_fpga_rdata_axi_s1_i95                =>  fabric_fpga_rdata_axi_s1_i(94)
       , fabric_fpga_rdata_axi_s1_i96                =>  fabric_fpga_rdata_axi_s1_i(95)
       , fabric_fpga_rdata_axi_s1_i97                =>  fabric_fpga_rdata_axi_s1_i(96)
       , fabric_fpga_rdata_axi_s1_i98                =>  fabric_fpga_rdata_axi_s1_i(97)
       , fabric_fpga_rdata_axi_s1_i99                =>  fabric_fpga_rdata_axi_s1_i(98)
       , fabric_fpga_rdata_axi_s1_i100               =>  fabric_fpga_rdata_axi_s1_i(99)
       , fabric_fpga_rdata_axi_s1_i101               =>  fabric_fpga_rdata_axi_s1_i(100)
       , fabric_fpga_rdata_axi_s1_i102               =>  fabric_fpga_rdata_axi_s1_i(101)
       , fabric_fpga_rdata_axi_s1_i103               =>  fabric_fpga_rdata_axi_s1_i(102)
       , fabric_fpga_rdata_axi_s1_i104               =>  fabric_fpga_rdata_axi_s1_i(103)
       , fabric_fpga_rdata_axi_s1_i105               =>  fabric_fpga_rdata_axi_s1_i(104)
       , fabric_fpga_rdata_axi_s1_i106               =>  fabric_fpga_rdata_axi_s1_i(105)
       , fabric_fpga_rdata_axi_s1_i107               =>  fabric_fpga_rdata_axi_s1_i(106)
       , fabric_fpga_rdata_axi_s1_i108               =>  fabric_fpga_rdata_axi_s1_i(107)
       , fabric_fpga_rdata_axi_s1_i109               =>  fabric_fpga_rdata_axi_s1_i(108)
       , fabric_fpga_rdata_axi_s1_i110               =>  fabric_fpga_rdata_axi_s1_i(109)
       , fabric_fpga_rdata_axi_s1_i111               =>  fabric_fpga_rdata_axi_s1_i(110)
       , fabric_fpga_rdata_axi_s1_i112               =>  fabric_fpga_rdata_axi_s1_i(111)
       , fabric_fpga_rdata_axi_s1_i113               =>  fabric_fpga_rdata_axi_s1_i(112)
       , fabric_fpga_rdata_axi_s1_i114               =>  fabric_fpga_rdata_axi_s1_i(113)
       , fabric_fpga_rdata_axi_s1_i115               =>  fabric_fpga_rdata_axi_s1_i(114)
       , fabric_fpga_rdata_axi_s1_i116               =>  fabric_fpga_rdata_axi_s1_i(115)
       , fabric_fpga_rdata_axi_s1_i117               =>  fabric_fpga_rdata_axi_s1_i(116)
       , fabric_fpga_rdata_axi_s1_i118               =>  fabric_fpga_rdata_axi_s1_i(117)
       , fabric_fpga_rdata_axi_s1_i119               =>  fabric_fpga_rdata_axi_s1_i(118)
       , fabric_fpga_rdata_axi_s1_i120               =>  fabric_fpga_rdata_axi_s1_i(119)
       , fabric_fpga_rdata_axi_s1_i121               =>  fabric_fpga_rdata_axi_s1_i(120)
       , fabric_fpga_rdata_axi_s1_i122               =>  fabric_fpga_rdata_axi_s1_i(121)
       , fabric_fpga_rdata_axi_s1_i123               =>  fabric_fpga_rdata_axi_s1_i(122)
       , fabric_fpga_rdata_axi_s1_i124               =>  fabric_fpga_rdata_axi_s1_i(123)
       , fabric_fpga_rdata_axi_s1_i125               =>  fabric_fpga_rdata_axi_s1_i(124)
       , fabric_fpga_rdata_axi_s1_i126               =>  fabric_fpga_rdata_axi_s1_i(125)
       , fabric_fpga_rdata_axi_s1_i127               =>  fabric_fpga_rdata_axi_s1_i(126)
       , fabric_fpga_rdata_axi_s1_i128               =>  fabric_fpga_rdata_axi_s1_i(127)
       , fabric_fpga_rid_axi_s1_i1                   =>  fabric_fpga_rid_axi_s1_i(0)
       , fabric_fpga_rid_axi_s1_i2                   =>  fabric_fpga_rid_axi_s1_i(1)
       , fabric_fpga_rid_axi_s1_i3                   =>  fabric_fpga_rid_axi_s1_i(2)
       , fabric_fpga_rid_axi_s1_i4                   =>  fabric_fpga_rid_axi_s1_i(3)
       , fabric_fpga_rid_axi_s1_i5                   =>  fabric_fpga_rid_axi_s1_i(4)
       , fabric_fpga_rid_axi_s1_i6                   =>  fabric_fpga_rid_axi_s1_i(5)
       , fabric_fpga_rid_axi_s1_i7                   =>  fabric_fpga_rid_axi_s1_i(6)
       , fabric_fpga_rid_axi_s1_i8                   =>  fabric_fpga_rid_axi_s1_i(7)
       , fabric_fpga_rid_axi_s1_i9                   =>  fabric_fpga_rid_axi_s1_i(8)
       , fabric_fpga_rid_axi_s1_i10                  =>  fabric_fpga_rid_axi_s1_i(9)
       , fabric_fpga_rid_axi_s1_i11                  =>  fabric_fpga_rid_axi_s1_i(10)
       , fabric_fpga_rid_axi_s1_i12                  =>  fabric_fpga_rid_axi_s1_i(11)
       , fabric_fpga_rlast_axi_s1_i                  =>  fabric_fpga_rlast_axi_s1_i
       , fabric_fpga_rresp_axi_s1_i1                 =>  fabric_fpga_rresp_axi_s1_i(0)
       , fabric_fpga_rresp_axi_s1_i2                 =>  fabric_fpga_rresp_axi_s1_i(1)
       , fabric_fpga_rvalid_axi_s1_i                 =>  fabric_fpga_rvalid_axi_s1_i
       , fabric_fpga_wready_axi_s1_i                 =>  fabric_fpga_wready_axi_s1_i
       , fabric_fpga_araddr_axi_s2_o1                =>  fabric_fpga_araddr_axi_s2_o(0)
       , fabric_fpga_araddr_axi_s2_o2                =>  fabric_fpga_araddr_axi_s2_o(1)
       , fabric_fpga_araddr_axi_s2_o3                =>  fabric_fpga_araddr_axi_s2_o(2)
       , fabric_fpga_araddr_axi_s2_o4                =>  fabric_fpga_araddr_axi_s2_o(3)
       , fabric_fpga_araddr_axi_s2_o5                =>  fabric_fpga_araddr_axi_s2_o(4)
       , fabric_fpga_araddr_axi_s2_o6                =>  fabric_fpga_araddr_axi_s2_o(5)
       , fabric_fpga_araddr_axi_s2_o7                =>  fabric_fpga_araddr_axi_s2_o(6)
       , fabric_fpga_araddr_axi_s2_o8                =>  fabric_fpga_araddr_axi_s2_o(7)
       , fabric_fpga_araddr_axi_s2_o9                =>  fabric_fpga_araddr_axi_s2_o(8)
       , fabric_fpga_araddr_axi_s2_o10               =>  fabric_fpga_araddr_axi_s2_o(9)
       , fabric_fpga_araddr_axi_s2_o11               =>  fabric_fpga_araddr_axi_s2_o(10)
       , fabric_fpga_araddr_axi_s2_o12               =>  fabric_fpga_araddr_axi_s2_o(11)
       , fabric_fpga_araddr_axi_s2_o13               =>  fabric_fpga_araddr_axi_s2_o(12)
       , fabric_fpga_araddr_axi_s2_o14               =>  fabric_fpga_araddr_axi_s2_o(13)
       , fabric_fpga_araddr_axi_s2_o15               =>  fabric_fpga_araddr_axi_s2_o(14)
       , fabric_fpga_araddr_axi_s2_o16               =>  fabric_fpga_araddr_axi_s2_o(15)
       , fabric_fpga_araddr_axi_s2_o17               =>  fabric_fpga_araddr_axi_s2_o(16)
       , fabric_fpga_araddr_axi_s2_o18               =>  fabric_fpga_araddr_axi_s2_o(17)
       , fabric_fpga_araddr_axi_s2_o19               =>  fabric_fpga_araddr_axi_s2_o(18)
       , fabric_fpga_araddr_axi_s2_o20               =>  fabric_fpga_araddr_axi_s2_o(19)
       , fabric_fpga_araddr_axi_s2_o21               =>  fabric_fpga_araddr_axi_s2_o(20)
       , fabric_fpga_araddr_axi_s2_o22               =>  fabric_fpga_araddr_axi_s2_o(21)
       , fabric_fpga_araddr_axi_s2_o23               =>  fabric_fpga_araddr_axi_s2_o(22)
       , fabric_fpga_araddr_axi_s2_o24               =>  fabric_fpga_araddr_axi_s2_o(23)
       , fabric_fpga_araddr_axi_s2_o25               =>  fabric_fpga_araddr_axi_s2_o(24)
       , fabric_fpga_araddr_axi_s2_o26               =>  fabric_fpga_araddr_axi_s2_o(25)
       , fabric_fpga_araddr_axi_s2_o27               =>  fabric_fpga_araddr_axi_s2_o(26)
       , fabric_fpga_araddr_axi_s2_o28               =>  fabric_fpga_araddr_axi_s2_o(27)
       , fabric_fpga_araddr_axi_s2_o29               =>  fabric_fpga_araddr_axi_s2_o(28)
       , fabric_fpga_araddr_axi_s2_o30               =>  fabric_fpga_araddr_axi_s2_o(29)
       , fabric_fpga_araddr_axi_s2_o31               =>  fabric_fpga_araddr_axi_s2_o(30)
       , fabric_fpga_araddr_axi_s2_o32               =>  fabric_fpga_araddr_axi_s2_o(31)
       , fabric_fpga_araddr_axi_s2_o33               =>  fabric_fpga_araddr_axi_s2_o(32)
       , fabric_fpga_araddr_axi_s2_o34               =>  fabric_fpga_araddr_axi_s2_o(33)
       , fabric_fpga_araddr_axi_s2_o35               =>  fabric_fpga_araddr_axi_s2_o(34)
       , fabric_fpga_araddr_axi_s2_o36               =>  fabric_fpga_araddr_axi_s2_o(35)
       , fabric_fpga_araddr_axi_s2_o37               =>  fabric_fpga_araddr_axi_s2_o(36)
       , fabric_fpga_araddr_axi_s2_o38               =>  fabric_fpga_araddr_axi_s2_o(37)
       , fabric_fpga_araddr_axi_s2_o39               =>  fabric_fpga_araddr_axi_s2_o(38)
       , fabric_fpga_araddr_axi_s2_o40               =>  fabric_fpga_araddr_axi_s2_o(39)
       , fabric_fpga_arburst_axi_s2_o1               =>  fabric_fpga_arburst_axi_s2_o(0)
       , fabric_fpga_arburst_axi_s2_o2               =>  fabric_fpga_arburst_axi_s2_o(1)
       , fabric_fpga_arcache_axi_s2_o1               =>  fabric_fpga_arcache_axi_s2_o(0)
       , fabric_fpga_arcache_axi_s2_o2               =>  fabric_fpga_arcache_axi_s2_o(1)
       , fabric_fpga_arcache_axi_s2_o3               =>  fabric_fpga_arcache_axi_s2_o(2)
       , fabric_fpga_arcache_axi_s2_o4               =>  fabric_fpga_arcache_axi_s2_o(3)
       , fabric_fpga_arid_axi_s2_o1                  =>  fabric_fpga_arid_axi_s2_o(0)
       , fabric_fpga_arid_axi_s2_o2                  =>  fabric_fpga_arid_axi_s2_o(1)
       , fabric_fpga_arid_axi_s2_o3                  =>  fabric_fpga_arid_axi_s2_o(2)
       , fabric_fpga_arid_axi_s2_o4                  =>  fabric_fpga_arid_axi_s2_o(3)
       , fabric_fpga_arid_axi_s2_o5                  =>  fabric_fpga_arid_axi_s2_o(4)
       , fabric_fpga_arid_axi_s2_o6                  =>  fabric_fpga_arid_axi_s2_o(5)
       , fabric_fpga_arid_axi_s2_o7                  =>  fabric_fpga_arid_axi_s2_o(6)
       , fabric_fpga_arid_axi_s2_o8                  =>  fabric_fpga_arid_axi_s2_o(7)
       , fabric_fpga_arid_axi_s2_o9                  =>  fabric_fpga_arid_axi_s2_o(8)
       , fabric_fpga_arid_axi_s2_o10                 =>  fabric_fpga_arid_axi_s2_o(9)
       , fabric_fpga_arid_axi_s2_o11                 =>  fabric_fpga_arid_axi_s2_o(10)
       , fabric_fpga_arid_axi_s2_o12                 =>  fabric_fpga_arid_axi_s2_o(11)
       , fabric_fpga_arlen_axi_s2_o1                 =>  fabric_fpga_arlen_axi_s2_o(0)
       , fabric_fpga_arlen_axi_s2_o2                 =>  fabric_fpga_arlen_axi_s2_o(1)
       , fabric_fpga_arlen_axi_s2_o3                 =>  fabric_fpga_arlen_axi_s2_o(2)
       , fabric_fpga_arlen_axi_s2_o4                 =>  fabric_fpga_arlen_axi_s2_o(3)
       , fabric_fpga_arlen_axi_s2_o5                 =>  fabric_fpga_arlen_axi_s2_o(4)
       , fabric_fpga_arlen_axi_s2_o6                 =>  fabric_fpga_arlen_axi_s2_o(5)
       , fabric_fpga_arlen_axi_s2_o7                 =>  fabric_fpga_arlen_axi_s2_o(6)
       , fabric_fpga_arlen_axi_s2_o8                 =>  fabric_fpga_arlen_axi_s2_o(7)
       , fabric_fpga_arlock_axi_s2_o                 =>  fabric_fpga_arlock_axi_s2_o
       , fabric_fpga_arprot_axi_s2_o1                =>  fabric_fpga_arprot_axi_s2_o(0)
       , fabric_fpga_arprot_axi_s2_o2                =>  fabric_fpga_arprot_axi_s2_o(1)
       , fabric_fpga_arprot_axi_s2_o3                =>  fabric_fpga_arprot_axi_s2_o(2)
       , fabric_fpga_arqos_axi_s2_o1                 =>  fabric_fpga_arqos_axi_s2_o(0)
       , fabric_fpga_arqos_axi_s2_o2                 =>  fabric_fpga_arqos_axi_s2_o(1)
       , fabric_fpga_arqos_axi_s2_o3                 =>  fabric_fpga_arqos_axi_s2_o(2)
       , fabric_fpga_arqos_axi_s2_o4                 =>  fabric_fpga_arqos_axi_s2_o(3)
       , fabric_fpga_arregion_axi_s2_o1              =>  fabric_fpga_arregion_axi_s2_o(0)
       , fabric_fpga_arregion_axi_s2_o2              =>  fabric_fpga_arregion_axi_s2_o(1)
       , fabric_fpga_arregion_axi_s2_o3              =>  fabric_fpga_arregion_axi_s2_o(2)
       , fabric_fpga_arregion_axi_s2_o4              =>  fabric_fpga_arregion_axi_s2_o(3)
       , fabric_fpga_arsize_axi_s2_o1                =>  fabric_fpga_arsize_axi_s2_o(0)
       , fabric_fpga_arsize_axi_s2_o2                =>  fabric_fpga_arsize_axi_s2_o(1)
       , fabric_fpga_arsize_axi_s2_o3                =>  fabric_fpga_arsize_axi_s2_o(2)
       , fabric_fpga_arvalid_axi_s2_o                =>  fabric_fpga_arvalid_axi_s2_o
       , fabric_fpga_awaddr_axi_s2_o1                =>  fabric_fpga_awaddr_axi_s2_o(0)
       , fabric_fpga_awaddr_axi_s2_o2                =>  fabric_fpga_awaddr_axi_s2_o(1)
       , fabric_fpga_awaddr_axi_s2_o3                =>  fabric_fpga_awaddr_axi_s2_o(2)
       , fabric_fpga_awaddr_axi_s2_o4                =>  fabric_fpga_awaddr_axi_s2_o(3)
       , fabric_fpga_awaddr_axi_s2_o5                =>  fabric_fpga_awaddr_axi_s2_o(4)
       , fabric_fpga_awaddr_axi_s2_o6                =>  fabric_fpga_awaddr_axi_s2_o(5)
       , fabric_fpga_awaddr_axi_s2_o7                =>  fabric_fpga_awaddr_axi_s2_o(6)
       , fabric_fpga_awaddr_axi_s2_o8                =>  fabric_fpga_awaddr_axi_s2_o(7)
       , fabric_fpga_awaddr_axi_s2_o9                =>  fabric_fpga_awaddr_axi_s2_o(8)
       , fabric_fpga_awaddr_axi_s2_o10               =>  fabric_fpga_awaddr_axi_s2_o(9)
       , fabric_fpga_awaddr_axi_s2_o11               =>  fabric_fpga_awaddr_axi_s2_o(10)
       , fabric_fpga_awaddr_axi_s2_o12               =>  fabric_fpga_awaddr_axi_s2_o(11)
       , fabric_fpga_awaddr_axi_s2_o13               =>  fabric_fpga_awaddr_axi_s2_o(12)
       , fabric_fpga_awaddr_axi_s2_o14               =>  fabric_fpga_awaddr_axi_s2_o(13)
       , fabric_fpga_awaddr_axi_s2_o15               =>  fabric_fpga_awaddr_axi_s2_o(14)
       , fabric_fpga_awaddr_axi_s2_o16               =>  fabric_fpga_awaddr_axi_s2_o(15)
       , fabric_fpga_awaddr_axi_s2_o17               =>  fabric_fpga_awaddr_axi_s2_o(16)
       , fabric_fpga_awaddr_axi_s2_o18               =>  fabric_fpga_awaddr_axi_s2_o(17)
       , fabric_fpga_awaddr_axi_s2_o19               =>  fabric_fpga_awaddr_axi_s2_o(18)
       , fabric_fpga_awaddr_axi_s2_o20               =>  fabric_fpga_awaddr_axi_s2_o(19)
       , fabric_fpga_awaddr_axi_s2_o21               =>  fabric_fpga_awaddr_axi_s2_o(20)
       , fabric_fpga_awaddr_axi_s2_o22               =>  fabric_fpga_awaddr_axi_s2_o(21)
       , fabric_fpga_awaddr_axi_s2_o23               =>  fabric_fpga_awaddr_axi_s2_o(22)
       , fabric_fpga_awaddr_axi_s2_o24               =>  fabric_fpga_awaddr_axi_s2_o(23)
       , fabric_fpga_awaddr_axi_s2_o25               =>  fabric_fpga_awaddr_axi_s2_o(24)
       , fabric_fpga_awaddr_axi_s2_o26               =>  fabric_fpga_awaddr_axi_s2_o(25)
       , fabric_fpga_awaddr_axi_s2_o27               =>  fabric_fpga_awaddr_axi_s2_o(26)
       , fabric_fpga_awaddr_axi_s2_o28               =>  fabric_fpga_awaddr_axi_s2_o(27)
       , fabric_fpga_awaddr_axi_s2_o29               =>  fabric_fpga_awaddr_axi_s2_o(28)
       , fabric_fpga_awaddr_axi_s2_o30               =>  fabric_fpga_awaddr_axi_s2_o(29)
       , fabric_fpga_awaddr_axi_s2_o31               =>  fabric_fpga_awaddr_axi_s2_o(30)
       , fabric_fpga_awaddr_axi_s2_o32               =>  fabric_fpga_awaddr_axi_s2_o(31)
       , fabric_fpga_awaddr_axi_s2_o33               =>  fabric_fpga_awaddr_axi_s2_o(32)
       , fabric_fpga_awaddr_axi_s2_o34               =>  fabric_fpga_awaddr_axi_s2_o(33)
       , fabric_fpga_awaddr_axi_s2_o35               =>  fabric_fpga_awaddr_axi_s2_o(34)
       , fabric_fpga_awaddr_axi_s2_o36               =>  fabric_fpga_awaddr_axi_s2_o(35)
       , fabric_fpga_awaddr_axi_s2_o37               =>  fabric_fpga_awaddr_axi_s2_o(36)
       , fabric_fpga_awaddr_axi_s2_o38               =>  fabric_fpga_awaddr_axi_s2_o(37)
       , fabric_fpga_awaddr_axi_s2_o39               =>  fabric_fpga_awaddr_axi_s2_o(38)
       , fabric_fpga_awaddr_axi_s2_o40               =>  fabric_fpga_awaddr_axi_s2_o(39)
       , fabric_fpga_awburst_axi_s2_o1               =>  fabric_fpga_awburst_axi_s2_o(0)
       , fabric_fpga_awburst_axi_s2_o2               =>  fabric_fpga_awburst_axi_s2_o(1)
       , fabric_fpga_awcache_axi_s2_o1               =>  fabric_fpga_awcache_axi_s2_o(0)
       , fabric_fpga_awcache_axi_s2_o2               =>  fabric_fpga_awcache_axi_s2_o(1)
       , fabric_fpga_awcache_axi_s2_o3               =>  fabric_fpga_awcache_axi_s2_o(2)
       , fabric_fpga_awcache_axi_s2_o4               =>  fabric_fpga_awcache_axi_s2_o(3)
       , fabric_fpga_awid_axi_s2_o1                  =>  fabric_fpga_awid_axi_s2_o(0)
       , fabric_fpga_awid_axi_s2_o2                  =>  fabric_fpga_awid_axi_s2_o(1)
       , fabric_fpga_awid_axi_s2_o3                  =>  fabric_fpga_awid_axi_s2_o(2)
       , fabric_fpga_awid_axi_s2_o4                  =>  fabric_fpga_awid_axi_s2_o(3)
       , fabric_fpga_awid_axi_s2_o5                  =>  fabric_fpga_awid_axi_s2_o(4)
       , fabric_fpga_awid_axi_s2_o6                  =>  fabric_fpga_awid_axi_s2_o(5)
       , fabric_fpga_awid_axi_s2_o7                  =>  fabric_fpga_awid_axi_s2_o(6)
       , fabric_fpga_awid_axi_s2_o8                  =>  fabric_fpga_awid_axi_s2_o(7)
       , fabric_fpga_awid_axi_s2_o9                  =>  fabric_fpga_awid_axi_s2_o(8)
       , fabric_fpga_awid_axi_s2_o10                 =>  fabric_fpga_awid_axi_s2_o(9)
       , fabric_fpga_awid_axi_s2_o11                 =>  fabric_fpga_awid_axi_s2_o(10)
       , fabric_fpga_awid_axi_s2_o12                 =>  fabric_fpga_awid_axi_s2_o(11)
       , fabric_fpga_awlen_axi_s2_o1                 =>  fabric_fpga_awlen_axi_s2_o(0)
       , fabric_fpga_awlen_axi_s2_o2                 =>  fabric_fpga_awlen_axi_s2_o(1)
       , fabric_fpga_awlen_axi_s2_o3                 =>  fabric_fpga_awlen_axi_s2_o(2)
       , fabric_fpga_awlen_axi_s2_o4                 =>  fabric_fpga_awlen_axi_s2_o(3)
       , fabric_fpga_awlen_axi_s2_o5                 =>  fabric_fpga_awlen_axi_s2_o(4)
       , fabric_fpga_awlen_axi_s2_o6                 =>  fabric_fpga_awlen_axi_s2_o(5)
       , fabric_fpga_awlen_axi_s2_o7                 =>  fabric_fpga_awlen_axi_s2_o(6)
       , fabric_fpga_awlen_axi_s2_o8                 =>  fabric_fpga_awlen_axi_s2_o(7)
       , fabric_fpga_awlock_axi_s2_o                 =>  fabric_fpga_awlock_axi_s2_o
       , fabric_fpga_awprot_axi_s2_o1                =>  fabric_fpga_awprot_axi_s2_o(0)
       , fabric_fpga_awprot_axi_s2_o2                =>  fabric_fpga_awprot_axi_s2_o(1)
       , fabric_fpga_awprot_axi_s2_o3                =>  fabric_fpga_awprot_axi_s2_o(2)
       , fabric_fpga_awqos_axi_s2_o1                 =>  fabric_fpga_awqos_axi_s2_o(0)
       , fabric_fpga_awqos_axi_s2_o2                 =>  fabric_fpga_awqos_axi_s2_o(1)
       , fabric_fpga_awqos_axi_s2_o3                 =>  fabric_fpga_awqos_axi_s2_o(2)
       , fabric_fpga_awqos_axi_s2_o4                 =>  fabric_fpga_awqos_axi_s2_o(3)
       , fabric_fpga_awregion_axi_s2_o1              =>  fabric_fpga_awregion_axi_s2_o(0)
       , fabric_fpga_awregion_axi_s2_o2              =>  fabric_fpga_awregion_axi_s2_o(1)
       , fabric_fpga_awregion_axi_s2_o3              =>  fabric_fpga_awregion_axi_s2_o(2)
       , fabric_fpga_awregion_axi_s2_o4              =>  fabric_fpga_awregion_axi_s2_o(3)
       , fabric_fpga_awsize_axi_s2_o1                =>  fabric_fpga_awsize_axi_s2_o(0)
       , fabric_fpga_awsize_axi_s2_o2                =>  fabric_fpga_awsize_axi_s2_o(1)
       , fabric_fpga_awsize_axi_s2_o3                =>  fabric_fpga_awsize_axi_s2_o(2)
       , fabric_fpga_bready_axi_s2_o                 =>  fabric_fpga_bready_axi_s2_o
       , fabric_fpga_rready_axi_s2_o                 =>  fabric_fpga_rready_axi_s2_o
       , fabric_fpga_wdata_axi_s2_o1                 =>  fabric_fpga_wdata_axi_s2_o(0)
       , fabric_fpga_wdata_axi_s2_o2                 =>  fabric_fpga_wdata_axi_s2_o(1)
       , fabric_fpga_wdata_axi_s2_o3                 =>  fabric_fpga_wdata_axi_s2_o(2)
       , fabric_fpga_wdata_axi_s2_o4                 =>  fabric_fpga_wdata_axi_s2_o(3)
       , fabric_fpga_wdata_axi_s2_o5                 =>  fabric_fpga_wdata_axi_s2_o(4)
       , fabric_fpga_wdata_axi_s2_o6                 =>  fabric_fpga_wdata_axi_s2_o(5)
       , fabric_fpga_wdata_axi_s2_o7                 =>  fabric_fpga_wdata_axi_s2_o(6)
       , fabric_fpga_wdata_axi_s2_o8                 =>  fabric_fpga_wdata_axi_s2_o(7)
       , fabric_fpga_wdata_axi_s2_o9                 =>  fabric_fpga_wdata_axi_s2_o(8)
       , fabric_fpga_wdata_axi_s2_o10                =>  fabric_fpga_wdata_axi_s2_o(9)
       , fabric_fpga_wdata_axi_s2_o11                =>  fabric_fpga_wdata_axi_s2_o(10)
       , fabric_fpga_wdata_axi_s2_o12                =>  fabric_fpga_wdata_axi_s2_o(11)
       , fabric_fpga_wdata_axi_s2_o13                =>  fabric_fpga_wdata_axi_s2_o(12)
       , fabric_fpga_wdata_axi_s2_o14                =>  fabric_fpga_wdata_axi_s2_o(13)
       , fabric_fpga_wdata_axi_s2_o15                =>  fabric_fpga_wdata_axi_s2_o(14)
       , fabric_fpga_wdata_axi_s2_o16                =>  fabric_fpga_wdata_axi_s2_o(15)
       , fabric_fpga_wdata_axi_s2_o17                =>  fabric_fpga_wdata_axi_s2_o(16)
       , fabric_fpga_wdata_axi_s2_o18                =>  fabric_fpga_wdata_axi_s2_o(17)
       , fabric_fpga_wdata_axi_s2_o19                =>  fabric_fpga_wdata_axi_s2_o(18)
       , fabric_fpga_wdata_axi_s2_o20                =>  fabric_fpga_wdata_axi_s2_o(19)
       , fabric_fpga_wdata_axi_s2_o21                =>  fabric_fpga_wdata_axi_s2_o(20)
       , fabric_fpga_wdata_axi_s2_o22                =>  fabric_fpga_wdata_axi_s2_o(21)
       , fabric_fpga_wdata_axi_s2_o23                =>  fabric_fpga_wdata_axi_s2_o(22)
       , fabric_fpga_wdata_axi_s2_o24                =>  fabric_fpga_wdata_axi_s2_o(23)
       , fabric_fpga_wdata_axi_s2_o25                =>  fabric_fpga_wdata_axi_s2_o(24)
       , fabric_fpga_wdata_axi_s2_o26                =>  fabric_fpga_wdata_axi_s2_o(25)
       , fabric_fpga_wdata_axi_s2_o27                =>  fabric_fpga_wdata_axi_s2_o(26)
       , fabric_fpga_wdata_axi_s2_o28                =>  fabric_fpga_wdata_axi_s2_o(27)
       , fabric_fpga_wdata_axi_s2_o29                =>  fabric_fpga_wdata_axi_s2_o(28)
       , fabric_fpga_wdata_axi_s2_o30                =>  fabric_fpga_wdata_axi_s2_o(29)
       , fabric_fpga_wdata_axi_s2_o31                =>  fabric_fpga_wdata_axi_s2_o(30)
       , fabric_fpga_wdata_axi_s2_o32                =>  fabric_fpga_wdata_axi_s2_o(31)
       , fabric_fpga_wdata_axi_s2_o33                =>  fabric_fpga_wdata_axi_s2_o(32)
       , fabric_fpga_wdata_axi_s2_o34                =>  fabric_fpga_wdata_axi_s2_o(33)
       , fabric_fpga_wdata_axi_s2_o35                =>  fabric_fpga_wdata_axi_s2_o(34)
       , fabric_fpga_wdata_axi_s2_o36                =>  fabric_fpga_wdata_axi_s2_o(35)
       , fabric_fpga_wdata_axi_s2_o37                =>  fabric_fpga_wdata_axi_s2_o(36)
       , fabric_fpga_wdata_axi_s2_o38                =>  fabric_fpga_wdata_axi_s2_o(37)
       , fabric_fpga_wdata_axi_s2_o39                =>  fabric_fpga_wdata_axi_s2_o(38)
       , fabric_fpga_wdata_axi_s2_o40                =>  fabric_fpga_wdata_axi_s2_o(39)
       , fabric_fpga_wdata_axi_s2_o41                =>  fabric_fpga_wdata_axi_s2_o(40)
       , fabric_fpga_wdata_axi_s2_o42                =>  fabric_fpga_wdata_axi_s2_o(41)
       , fabric_fpga_wdata_axi_s2_o43                =>  fabric_fpga_wdata_axi_s2_o(42)
       , fabric_fpga_wdata_axi_s2_o44                =>  fabric_fpga_wdata_axi_s2_o(43)
       , fabric_fpga_wdata_axi_s2_o45                =>  fabric_fpga_wdata_axi_s2_o(44)
       , fabric_fpga_wdata_axi_s2_o46                =>  fabric_fpga_wdata_axi_s2_o(45)
       , fabric_fpga_wdata_axi_s2_o47                =>  fabric_fpga_wdata_axi_s2_o(46)
       , fabric_fpga_wdata_axi_s2_o48                =>  fabric_fpga_wdata_axi_s2_o(47)
       , fabric_fpga_wdata_axi_s2_o49                =>  fabric_fpga_wdata_axi_s2_o(48)
       , fabric_fpga_wdata_axi_s2_o50                =>  fabric_fpga_wdata_axi_s2_o(49)
       , fabric_fpga_wdata_axi_s2_o51                =>  fabric_fpga_wdata_axi_s2_o(50)
       , fabric_fpga_wdata_axi_s2_o52                =>  fabric_fpga_wdata_axi_s2_o(51)
       , fabric_fpga_wdata_axi_s2_o53                =>  fabric_fpga_wdata_axi_s2_o(52)
       , fabric_fpga_wdata_axi_s2_o54                =>  fabric_fpga_wdata_axi_s2_o(53)
       , fabric_fpga_wdata_axi_s2_o55                =>  fabric_fpga_wdata_axi_s2_o(54)
       , fabric_fpga_wdata_axi_s2_o56                =>  fabric_fpga_wdata_axi_s2_o(55)
       , fabric_fpga_wdata_axi_s2_o57                =>  fabric_fpga_wdata_axi_s2_o(56)
       , fabric_fpga_wdata_axi_s2_o58                =>  fabric_fpga_wdata_axi_s2_o(57)
       , fabric_fpga_wdata_axi_s2_o59                =>  fabric_fpga_wdata_axi_s2_o(58)
       , fabric_fpga_wdata_axi_s2_o60                =>  fabric_fpga_wdata_axi_s2_o(59)
       , fabric_fpga_wdata_axi_s2_o61                =>  fabric_fpga_wdata_axi_s2_o(60)
       , fabric_fpga_wdata_axi_s2_o62                =>  fabric_fpga_wdata_axi_s2_o(61)
       , fabric_fpga_wdata_axi_s2_o63                =>  fabric_fpga_wdata_axi_s2_o(62)
       , fabric_fpga_wdata_axi_s2_o64                =>  fabric_fpga_wdata_axi_s2_o(63)
       , fabric_fpga_wdata_axi_s2_o65                =>  fabric_fpga_wdata_axi_s2_o(64)
       , fabric_fpga_wdata_axi_s2_o66                =>  fabric_fpga_wdata_axi_s2_o(65)
       , fabric_fpga_wdata_axi_s2_o67                =>  fabric_fpga_wdata_axi_s2_o(66)
       , fabric_fpga_wdata_axi_s2_o68                =>  fabric_fpga_wdata_axi_s2_o(67)
       , fabric_fpga_wdata_axi_s2_o69                =>  fabric_fpga_wdata_axi_s2_o(68)
       , fabric_fpga_wdata_axi_s2_o70                =>  fabric_fpga_wdata_axi_s2_o(69)
       , fabric_fpga_wdata_axi_s2_o71                =>  fabric_fpga_wdata_axi_s2_o(70)
       , fabric_fpga_wdata_axi_s2_o72                =>  fabric_fpga_wdata_axi_s2_o(71)
       , fabric_fpga_wdata_axi_s2_o73                =>  fabric_fpga_wdata_axi_s2_o(72)
       , fabric_fpga_wdata_axi_s2_o74                =>  fabric_fpga_wdata_axi_s2_o(73)
       , fabric_fpga_wdata_axi_s2_o75                =>  fabric_fpga_wdata_axi_s2_o(74)
       , fabric_fpga_wdata_axi_s2_o76                =>  fabric_fpga_wdata_axi_s2_o(75)
       , fabric_fpga_wdata_axi_s2_o77                =>  fabric_fpga_wdata_axi_s2_o(76)
       , fabric_fpga_wdata_axi_s2_o78                =>  fabric_fpga_wdata_axi_s2_o(77)
       , fabric_fpga_wdata_axi_s2_o79                =>  fabric_fpga_wdata_axi_s2_o(78)
       , fabric_fpga_wdata_axi_s2_o80                =>  fabric_fpga_wdata_axi_s2_o(79)
       , fabric_fpga_wdata_axi_s2_o81                =>  fabric_fpga_wdata_axi_s2_o(80)
       , fabric_fpga_wdata_axi_s2_o82                =>  fabric_fpga_wdata_axi_s2_o(81)
       , fabric_fpga_wdata_axi_s2_o83                =>  fabric_fpga_wdata_axi_s2_o(82)
       , fabric_fpga_wdata_axi_s2_o84                =>  fabric_fpga_wdata_axi_s2_o(83)
       , fabric_fpga_wdata_axi_s2_o85                =>  fabric_fpga_wdata_axi_s2_o(84)
       , fabric_fpga_wdata_axi_s2_o86                =>  fabric_fpga_wdata_axi_s2_o(85)
       , fabric_fpga_wdata_axi_s2_o87                =>  fabric_fpga_wdata_axi_s2_o(86)
       , fabric_fpga_wdata_axi_s2_o88                =>  fabric_fpga_wdata_axi_s2_o(87)
       , fabric_fpga_wdata_axi_s2_o89                =>  fabric_fpga_wdata_axi_s2_o(88)
       , fabric_fpga_wdata_axi_s2_o90                =>  fabric_fpga_wdata_axi_s2_o(89)
       , fabric_fpga_wdata_axi_s2_o91                =>  fabric_fpga_wdata_axi_s2_o(90)
       , fabric_fpga_wdata_axi_s2_o92                =>  fabric_fpga_wdata_axi_s2_o(91)
       , fabric_fpga_wdata_axi_s2_o93                =>  fabric_fpga_wdata_axi_s2_o(92)
       , fabric_fpga_wdata_axi_s2_o94                =>  fabric_fpga_wdata_axi_s2_o(93)
       , fabric_fpga_wdata_axi_s2_o95                =>  fabric_fpga_wdata_axi_s2_o(94)
       , fabric_fpga_wdata_axi_s2_o96                =>  fabric_fpga_wdata_axi_s2_o(95)
       , fabric_fpga_wdata_axi_s2_o97                =>  fabric_fpga_wdata_axi_s2_o(96)
       , fabric_fpga_wdata_axi_s2_o98                =>  fabric_fpga_wdata_axi_s2_o(97)
       , fabric_fpga_wdata_axi_s2_o99                =>  fabric_fpga_wdata_axi_s2_o(98)
       , fabric_fpga_wdata_axi_s2_o100               =>  fabric_fpga_wdata_axi_s2_o(99)
       , fabric_fpga_wdata_axi_s2_o101               =>  fabric_fpga_wdata_axi_s2_o(100)
       , fabric_fpga_wdata_axi_s2_o102               =>  fabric_fpga_wdata_axi_s2_o(101)
       , fabric_fpga_wdata_axi_s2_o103               =>  fabric_fpga_wdata_axi_s2_o(102)
       , fabric_fpga_wdata_axi_s2_o104               =>  fabric_fpga_wdata_axi_s2_o(103)
       , fabric_fpga_wdata_axi_s2_o105               =>  fabric_fpga_wdata_axi_s2_o(104)
       , fabric_fpga_wdata_axi_s2_o106               =>  fabric_fpga_wdata_axi_s2_o(105)
       , fabric_fpga_wdata_axi_s2_o107               =>  fabric_fpga_wdata_axi_s2_o(106)
       , fabric_fpga_wdata_axi_s2_o108               =>  fabric_fpga_wdata_axi_s2_o(107)
       , fabric_fpga_wdata_axi_s2_o109               =>  fabric_fpga_wdata_axi_s2_o(108)
       , fabric_fpga_wdata_axi_s2_o110               =>  fabric_fpga_wdata_axi_s2_o(109)
       , fabric_fpga_wdata_axi_s2_o111               =>  fabric_fpga_wdata_axi_s2_o(110)
       , fabric_fpga_wdata_axi_s2_o112               =>  fabric_fpga_wdata_axi_s2_o(111)
       , fabric_fpga_wdata_axi_s2_o113               =>  fabric_fpga_wdata_axi_s2_o(112)
       , fabric_fpga_wdata_axi_s2_o114               =>  fabric_fpga_wdata_axi_s2_o(113)
       , fabric_fpga_wdata_axi_s2_o115               =>  fabric_fpga_wdata_axi_s2_o(114)
       , fabric_fpga_wdata_axi_s2_o116               =>  fabric_fpga_wdata_axi_s2_o(115)
       , fabric_fpga_wdata_axi_s2_o117               =>  fabric_fpga_wdata_axi_s2_o(116)
       , fabric_fpga_wdata_axi_s2_o118               =>  fabric_fpga_wdata_axi_s2_o(117)
       , fabric_fpga_wdata_axi_s2_o119               =>  fabric_fpga_wdata_axi_s2_o(118)
       , fabric_fpga_wdata_axi_s2_o120               =>  fabric_fpga_wdata_axi_s2_o(119)
       , fabric_fpga_wdata_axi_s2_o121               =>  fabric_fpga_wdata_axi_s2_o(120)
       , fabric_fpga_wdata_axi_s2_o122               =>  fabric_fpga_wdata_axi_s2_o(121)
       , fabric_fpga_wdata_axi_s2_o123               =>  fabric_fpga_wdata_axi_s2_o(122)
       , fabric_fpga_wdata_axi_s2_o124               =>  fabric_fpga_wdata_axi_s2_o(123)
       , fabric_fpga_wdata_axi_s2_o125               =>  fabric_fpga_wdata_axi_s2_o(124)
       , fabric_fpga_wdata_axi_s2_o126               =>  fabric_fpga_wdata_axi_s2_o(125)
       , fabric_fpga_wdata_axi_s2_o127               =>  fabric_fpga_wdata_axi_s2_o(126)
       , fabric_fpga_wdata_axi_s2_o128               =>  fabric_fpga_wdata_axi_s2_o(127)
       , fabric_fpga_wlast_axi_s2_o                  =>  fabric_fpga_wlast_axi_s2_o
       , fabric_fpga_wstrb_axi_s2_o1                 =>  fabric_fpga_wstrb_axi_s2_o(0)
       , fabric_fpga_wstrb_axi_s2_o2                 =>  fabric_fpga_wstrb_axi_s2_o(1)
       , fabric_fpga_wstrb_axi_s2_o3                 =>  fabric_fpga_wstrb_axi_s2_o(2)
       , fabric_fpga_wstrb_axi_s2_o4                 =>  fabric_fpga_wstrb_axi_s2_o(3)
       , fabric_fpga_wstrb_axi_s2_o5                 =>  fabric_fpga_wstrb_axi_s2_o(4)
       , fabric_fpga_wstrb_axi_s2_o6                 =>  fabric_fpga_wstrb_axi_s2_o(5)
       , fabric_fpga_wstrb_axi_s2_o7                 =>  fabric_fpga_wstrb_axi_s2_o(6)
       , fabric_fpga_wstrb_axi_s2_o8                 =>  fabric_fpga_wstrb_axi_s2_o(7)
       , fabric_fpga_wstrb_axi_s2_o9                 =>  fabric_fpga_wstrb_axi_s2_o(8)
       , fabric_fpga_wstrb_axi_s2_o10                =>  fabric_fpga_wstrb_axi_s2_o(9)
       , fabric_fpga_wstrb_axi_s2_o11                =>  fabric_fpga_wstrb_axi_s2_o(10)
       , fabric_fpga_wstrb_axi_s2_o12                =>  fabric_fpga_wstrb_axi_s2_o(11)
       , fabric_fpga_wstrb_axi_s2_o13                =>  fabric_fpga_wstrb_axi_s2_o(12)
       , fabric_fpga_wstrb_axi_s2_o14                =>  fabric_fpga_wstrb_axi_s2_o(13)
       , fabric_fpga_wstrb_axi_s2_o15                =>  fabric_fpga_wstrb_axi_s2_o(14)
       , fabric_fpga_wstrb_axi_s2_o16                =>  fabric_fpga_wstrb_axi_s2_o(15)
       , fabric_fpga_wvalid_axi_s2_o                 =>  fabric_fpga_wvalid_axi_s2_o
       , fabric_fpga_awvalid_axi_s2_o                =>  fabric_fpga_awvalid_axi_s2_o
       , fabric_fpga_arready_axi_s2_i                =>  fabric_fpga_arready_axi_s2_i
       , fabric_fpga_awready_axi_s2_i                =>  fabric_fpga_awready_axi_s2_i
       , fabric_fpga_bid_axi_s2_i1                   =>  fabric_fpga_bid_axi_s2_i(0)
       , fabric_fpga_bid_axi_s2_i2                   =>  fabric_fpga_bid_axi_s2_i(1)
       , fabric_fpga_bid_axi_s2_i3                   =>  fabric_fpga_bid_axi_s2_i(2)
       , fabric_fpga_bid_axi_s2_i4                   =>  fabric_fpga_bid_axi_s2_i(3)
       , fabric_fpga_bid_axi_s2_i5                   =>  fabric_fpga_bid_axi_s2_i(4)
       , fabric_fpga_bid_axi_s2_i6                   =>  fabric_fpga_bid_axi_s2_i(5)
       , fabric_fpga_bid_axi_s2_i7                   =>  fabric_fpga_bid_axi_s2_i(6)
       , fabric_fpga_bid_axi_s2_i8                   =>  fabric_fpga_bid_axi_s2_i(7)
       , fabric_fpga_bid_axi_s2_i9                   =>  fabric_fpga_bid_axi_s2_i(8)
       , fabric_fpga_bid_axi_s2_i10                  =>  fabric_fpga_bid_axi_s2_i(9)
       , fabric_fpga_bid_axi_s2_i11                  =>  fabric_fpga_bid_axi_s2_i(10)
       , fabric_fpga_bid_axi_s2_i12                  =>  fabric_fpga_bid_axi_s2_i(11)
       , fabric_fpga_bresp_axi_s2_i1                 =>  fabric_fpga_bresp_axi_s2_i(0)
       , fabric_fpga_bresp_axi_s2_i2                 =>  fabric_fpga_bresp_axi_s2_i(1)
       , fabric_fpga_bvalid_axi_s2_i                 =>  fabric_fpga_bvalid_axi_s2_i
       , fabric_fpga_rdata_axi_s2_i1                 =>  fabric_fpga_rdata_axi_s2_i(0)
       , fabric_fpga_rdata_axi_s2_i2                 =>  fabric_fpga_rdata_axi_s2_i(1)
       , fabric_fpga_rdata_axi_s2_i3                 =>  fabric_fpga_rdata_axi_s2_i(2)
       , fabric_fpga_rdata_axi_s2_i4                 =>  fabric_fpga_rdata_axi_s2_i(3)
       , fabric_fpga_rdata_axi_s2_i5                 =>  fabric_fpga_rdata_axi_s2_i(4)
       , fabric_fpga_rdata_axi_s2_i6                 =>  fabric_fpga_rdata_axi_s2_i(5)
       , fabric_fpga_rdata_axi_s2_i7                 =>  fabric_fpga_rdata_axi_s2_i(6)
       , fabric_fpga_rdata_axi_s2_i8                 =>  fabric_fpga_rdata_axi_s2_i(7)
       , fabric_fpga_rdata_axi_s2_i9                 =>  fabric_fpga_rdata_axi_s2_i(8)
       , fabric_fpga_rdata_axi_s2_i10                =>  fabric_fpga_rdata_axi_s2_i(9)
       , fabric_fpga_rdata_axi_s2_i11                =>  fabric_fpga_rdata_axi_s2_i(10)
       , fabric_fpga_rdata_axi_s2_i12                =>  fabric_fpga_rdata_axi_s2_i(11)
       , fabric_fpga_rdata_axi_s2_i13                =>  fabric_fpga_rdata_axi_s2_i(12)
       , fabric_fpga_rdata_axi_s2_i14                =>  fabric_fpga_rdata_axi_s2_i(13)
       , fabric_fpga_rdata_axi_s2_i15                =>  fabric_fpga_rdata_axi_s2_i(14)
       , fabric_fpga_rdata_axi_s2_i16                =>  fabric_fpga_rdata_axi_s2_i(15)
       , fabric_fpga_rdata_axi_s2_i17                =>  fabric_fpga_rdata_axi_s2_i(16)
       , fabric_fpga_rdata_axi_s2_i18                =>  fabric_fpga_rdata_axi_s2_i(17)
       , fabric_fpga_rdata_axi_s2_i19                =>  fabric_fpga_rdata_axi_s2_i(18)
       , fabric_fpga_rdata_axi_s2_i20                =>  fabric_fpga_rdata_axi_s2_i(19)
       , fabric_fpga_rdata_axi_s2_i21                =>  fabric_fpga_rdata_axi_s2_i(20)
       , fabric_fpga_rdata_axi_s2_i22                =>  fabric_fpga_rdata_axi_s2_i(21)
       , fabric_fpga_rdata_axi_s2_i23                =>  fabric_fpga_rdata_axi_s2_i(22)
       , fabric_fpga_rdata_axi_s2_i24                =>  fabric_fpga_rdata_axi_s2_i(23)
       , fabric_fpga_rdata_axi_s2_i25                =>  fabric_fpga_rdata_axi_s2_i(24)
       , fabric_fpga_rdata_axi_s2_i26                =>  fabric_fpga_rdata_axi_s2_i(25)
       , fabric_fpga_rdata_axi_s2_i27                =>  fabric_fpga_rdata_axi_s2_i(26)
       , fabric_fpga_rdata_axi_s2_i28                =>  fabric_fpga_rdata_axi_s2_i(27)
       , fabric_fpga_rdata_axi_s2_i29                =>  fabric_fpga_rdata_axi_s2_i(28)
       , fabric_fpga_rdata_axi_s2_i30                =>  fabric_fpga_rdata_axi_s2_i(29)
       , fabric_fpga_rdata_axi_s2_i31                =>  fabric_fpga_rdata_axi_s2_i(30)
       , fabric_fpga_rdata_axi_s2_i32                =>  fabric_fpga_rdata_axi_s2_i(31)
       , fabric_fpga_rdata_axi_s2_i33                =>  fabric_fpga_rdata_axi_s2_i(32)
       , fabric_fpga_rdata_axi_s2_i34                =>  fabric_fpga_rdata_axi_s2_i(33)
       , fabric_fpga_rdata_axi_s2_i35                =>  fabric_fpga_rdata_axi_s2_i(34)
       , fabric_fpga_rdata_axi_s2_i36                =>  fabric_fpga_rdata_axi_s2_i(35)
       , fabric_fpga_rdata_axi_s2_i37                =>  fabric_fpga_rdata_axi_s2_i(36)
       , fabric_fpga_rdata_axi_s2_i38                =>  fabric_fpga_rdata_axi_s2_i(37)
       , fabric_fpga_rdata_axi_s2_i39                =>  fabric_fpga_rdata_axi_s2_i(38)
       , fabric_fpga_rdata_axi_s2_i40                =>  fabric_fpga_rdata_axi_s2_i(39)
       , fabric_fpga_rdata_axi_s2_i41                =>  fabric_fpga_rdata_axi_s2_i(40)
       , fabric_fpga_rdata_axi_s2_i42                =>  fabric_fpga_rdata_axi_s2_i(41)
       , fabric_fpga_rdata_axi_s2_i43                =>  fabric_fpga_rdata_axi_s2_i(42)
       , fabric_fpga_rdata_axi_s2_i44                =>  fabric_fpga_rdata_axi_s2_i(43)
       , fabric_fpga_rdata_axi_s2_i45                =>  fabric_fpga_rdata_axi_s2_i(44)
       , fabric_fpga_rdata_axi_s2_i46                =>  fabric_fpga_rdata_axi_s2_i(45)
       , fabric_fpga_rdata_axi_s2_i47                =>  fabric_fpga_rdata_axi_s2_i(46)
       , fabric_fpga_rdata_axi_s2_i48                =>  fabric_fpga_rdata_axi_s2_i(47)
       , fabric_fpga_rdata_axi_s2_i49                =>  fabric_fpga_rdata_axi_s2_i(48)
       , fabric_fpga_rdata_axi_s2_i50                =>  fabric_fpga_rdata_axi_s2_i(49)
       , fabric_fpga_rdata_axi_s2_i51                =>  fabric_fpga_rdata_axi_s2_i(50)
       , fabric_fpga_rdata_axi_s2_i52                =>  fabric_fpga_rdata_axi_s2_i(51)
       , fabric_fpga_rdata_axi_s2_i53                =>  fabric_fpga_rdata_axi_s2_i(52)
       , fabric_fpga_rdata_axi_s2_i54                =>  fabric_fpga_rdata_axi_s2_i(53)
       , fabric_fpga_rdata_axi_s2_i55                =>  fabric_fpga_rdata_axi_s2_i(54)
       , fabric_fpga_rdata_axi_s2_i56                =>  fabric_fpga_rdata_axi_s2_i(55)
       , fabric_fpga_rdata_axi_s2_i57                =>  fabric_fpga_rdata_axi_s2_i(56)
       , fabric_fpga_rdata_axi_s2_i58                =>  fabric_fpga_rdata_axi_s2_i(57)
       , fabric_fpga_rdata_axi_s2_i59                =>  fabric_fpga_rdata_axi_s2_i(58)
       , fabric_fpga_rdata_axi_s2_i60                =>  fabric_fpga_rdata_axi_s2_i(59)
       , fabric_fpga_rdata_axi_s2_i61                =>  fabric_fpga_rdata_axi_s2_i(60)
       , fabric_fpga_rdata_axi_s2_i62                =>  fabric_fpga_rdata_axi_s2_i(61)
       , fabric_fpga_rdata_axi_s2_i63                =>  fabric_fpga_rdata_axi_s2_i(62)
       , fabric_fpga_rdata_axi_s2_i64                =>  fabric_fpga_rdata_axi_s2_i(63)
       , fabric_fpga_rdata_axi_s2_i65                =>  fabric_fpga_rdata_axi_s2_i(64)
       , fabric_fpga_rdata_axi_s2_i66                =>  fabric_fpga_rdata_axi_s2_i(65)
       , fabric_fpga_rdata_axi_s2_i67                =>  fabric_fpga_rdata_axi_s2_i(66)
       , fabric_fpga_rdata_axi_s2_i68                =>  fabric_fpga_rdata_axi_s2_i(67)
       , fabric_fpga_rdata_axi_s2_i69                =>  fabric_fpga_rdata_axi_s2_i(68)
       , fabric_fpga_rdata_axi_s2_i70                =>  fabric_fpga_rdata_axi_s2_i(69)
       , fabric_fpga_rdata_axi_s2_i71                =>  fabric_fpga_rdata_axi_s2_i(70)
       , fabric_fpga_rdata_axi_s2_i72                =>  fabric_fpga_rdata_axi_s2_i(71)
       , fabric_fpga_rdata_axi_s2_i73                =>  fabric_fpga_rdata_axi_s2_i(72)
       , fabric_fpga_rdata_axi_s2_i74                =>  fabric_fpga_rdata_axi_s2_i(73)
       , fabric_fpga_rdata_axi_s2_i75                =>  fabric_fpga_rdata_axi_s2_i(74)
       , fabric_fpga_rdata_axi_s2_i76                =>  fabric_fpga_rdata_axi_s2_i(75)
       , fabric_fpga_rdata_axi_s2_i77                =>  fabric_fpga_rdata_axi_s2_i(76)
       , fabric_fpga_rdata_axi_s2_i78                =>  fabric_fpga_rdata_axi_s2_i(77)
       , fabric_fpga_rdata_axi_s2_i79                =>  fabric_fpga_rdata_axi_s2_i(78)
       , fabric_fpga_rdata_axi_s2_i80                =>  fabric_fpga_rdata_axi_s2_i(79)
       , fabric_fpga_rdata_axi_s2_i81                =>  fabric_fpga_rdata_axi_s2_i(80)
       , fabric_fpga_rdata_axi_s2_i82                =>  fabric_fpga_rdata_axi_s2_i(81)
       , fabric_fpga_rdata_axi_s2_i83                =>  fabric_fpga_rdata_axi_s2_i(82)
       , fabric_fpga_rdata_axi_s2_i84                =>  fabric_fpga_rdata_axi_s2_i(83)
       , fabric_fpga_rdata_axi_s2_i85                =>  fabric_fpga_rdata_axi_s2_i(84)
       , fabric_fpga_rdata_axi_s2_i86                =>  fabric_fpga_rdata_axi_s2_i(85)
       , fabric_fpga_rdata_axi_s2_i87                =>  fabric_fpga_rdata_axi_s2_i(86)
       , fabric_fpga_rdata_axi_s2_i88                =>  fabric_fpga_rdata_axi_s2_i(87)
       , fabric_fpga_rdata_axi_s2_i89                =>  fabric_fpga_rdata_axi_s2_i(88)
       , fabric_fpga_rdata_axi_s2_i90                =>  fabric_fpga_rdata_axi_s2_i(89)
       , fabric_fpga_rdata_axi_s2_i91                =>  fabric_fpga_rdata_axi_s2_i(90)
       , fabric_fpga_rdata_axi_s2_i92                =>  fabric_fpga_rdata_axi_s2_i(91)
       , fabric_fpga_rdata_axi_s2_i93                =>  fabric_fpga_rdata_axi_s2_i(92)
       , fabric_fpga_rdata_axi_s2_i94                =>  fabric_fpga_rdata_axi_s2_i(93)
       , fabric_fpga_rdata_axi_s2_i95                =>  fabric_fpga_rdata_axi_s2_i(94)
       , fabric_fpga_rdata_axi_s2_i96                =>  fabric_fpga_rdata_axi_s2_i(95)
       , fabric_fpga_rdata_axi_s2_i97                =>  fabric_fpga_rdata_axi_s2_i(96)
       , fabric_fpga_rdata_axi_s2_i98                =>  fabric_fpga_rdata_axi_s2_i(97)
       , fabric_fpga_rdata_axi_s2_i99                =>  fabric_fpga_rdata_axi_s2_i(98)
       , fabric_fpga_rdata_axi_s2_i100               =>  fabric_fpga_rdata_axi_s2_i(99)
       , fabric_fpga_rdata_axi_s2_i101               =>  fabric_fpga_rdata_axi_s2_i(100)
       , fabric_fpga_rdata_axi_s2_i102               =>  fabric_fpga_rdata_axi_s2_i(101)
       , fabric_fpga_rdata_axi_s2_i103               =>  fabric_fpga_rdata_axi_s2_i(102)
       , fabric_fpga_rdata_axi_s2_i104               =>  fabric_fpga_rdata_axi_s2_i(103)
       , fabric_fpga_rdata_axi_s2_i105               =>  fabric_fpga_rdata_axi_s2_i(104)
       , fabric_fpga_rdata_axi_s2_i106               =>  fabric_fpga_rdata_axi_s2_i(105)
       , fabric_fpga_rdata_axi_s2_i107               =>  fabric_fpga_rdata_axi_s2_i(106)
       , fabric_fpga_rdata_axi_s2_i108               =>  fabric_fpga_rdata_axi_s2_i(107)
       , fabric_fpga_rdata_axi_s2_i109               =>  fabric_fpga_rdata_axi_s2_i(108)
       , fabric_fpga_rdata_axi_s2_i110               =>  fabric_fpga_rdata_axi_s2_i(109)
       , fabric_fpga_rdata_axi_s2_i111               =>  fabric_fpga_rdata_axi_s2_i(110)
       , fabric_fpga_rdata_axi_s2_i112               =>  fabric_fpga_rdata_axi_s2_i(111)
       , fabric_fpga_rdata_axi_s2_i113               =>  fabric_fpga_rdata_axi_s2_i(112)
       , fabric_fpga_rdata_axi_s2_i114               =>  fabric_fpga_rdata_axi_s2_i(113)
       , fabric_fpga_rdata_axi_s2_i115               =>  fabric_fpga_rdata_axi_s2_i(114)
       , fabric_fpga_rdata_axi_s2_i116               =>  fabric_fpga_rdata_axi_s2_i(115)
       , fabric_fpga_rdata_axi_s2_i117               =>  fabric_fpga_rdata_axi_s2_i(116)
       , fabric_fpga_rdata_axi_s2_i118               =>  fabric_fpga_rdata_axi_s2_i(117)
       , fabric_fpga_rdata_axi_s2_i119               =>  fabric_fpga_rdata_axi_s2_i(118)
       , fabric_fpga_rdata_axi_s2_i120               =>  fabric_fpga_rdata_axi_s2_i(119)
       , fabric_fpga_rdata_axi_s2_i121               =>  fabric_fpga_rdata_axi_s2_i(120)
       , fabric_fpga_rdata_axi_s2_i122               =>  fabric_fpga_rdata_axi_s2_i(121)
       , fabric_fpga_rdata_axi_s2_i123               =>  fabric_fpga_rdata_axi_s2_i(122)
       , fabric_fpga_rdata_axi_s2_i124               =>  fabric_fpga_rdata_axi_s2_i(123)
       , fabric_fpga_rdata_axi_s2_i125               =>  fabric_fpga_rdata_axi_s2_i(124)
       , fabric_fpga_rdata_axi_s2_i126               =>  fabric_fpga_rdata_axi_s2_i(125)
       , fabric_fpga_rdata_axi_s2_i127               =>  fabric_fpga_rdata_axi_s2_i(126)
       , fabric_fpga_rdata_axi_s2_i128               =>  fabric_fpga_rdata_axi_s2_i(127)
       , fabric_fpga_rid_axi_s2_i1                   =>  fabric_fpga_rid_axi_s2_i(0)
       , fabric_fpga_rid_axi_s2_i2                   =>  fabric_fpga_rid_axi_s2_i(1)
       , fabric_fpga_rid_axi_s2_i3                   =>  fabric_fpga_rid_axi_s2_i(2)
       , fabric_fpga_rid_axi_s2_i4                   =>  fabric_fpga_rid_axi_s2_i(3)
       , fabric_fpga_rid_axi_s2_i5                   =>  fabric_fpga_rid_axi_s2_i(4)
       , fabric_fpga_rid_axi_s2_i6                   =>  fabric_fpga_rid_axi_s2_i(5)
       , fabric_fpga_rid_axi_s2_i7                   =>  fabric_fpga_rid_axi_s2_i(6)
       , fabric_fpga_rid_axi_s2_i8                   =>  fabric_fpga_rid_axi_s2_i(7)
       , fabric_fpga_rid_axi_s2_i9                   =>  fabric_fpga_rid_axi_s2_i(8)
       , fabric_fpga_rid_axi_s2_i10                  =>  fabric_fpga_rid_axi_s2_i(9)
       , fabric_fpga_rid_axi_s2_i11                  =>  fabric_fpga_rid_axi_s2_i(10)
       , fabric_fpga_rid_axi_s2_i12                  =>  fabric_fpga_rid_axi_s2_i(11)
       , fabric_fpga_rlast_axi_s2_i                  =>  fabric_fpga_rlast_axi_s2_i
       , fabric_fpga_rresp_axi_s2_i1                 =>  fabric_fpga_rresp_axi_s2_i(0)
       , fabric_fpga_rresp_axi_s2_i2                 =>  fabric_fpga_rresp_axi_s2_i(1)
       , fabric_fpga_rvalid_axi_s2_i                 =>  fabric_fpga_rvalid_axi_s2_i
       , fabric_fpga_wready_axi_s2_i                 =>  fabric_fpga_wready_axi_s2_i
       , fabric_fpga_arready_axi_m1_o                =>  fabric_fpga_arready_axi_m1_o
       , fabric_fpga_awready_axi_m1_o                =>  fabric_fpga_awready_axi_m1_o
       , fabric_fpga_bid_axi_m1_o1                   =>  fabric_fpga_bid_axi_m1_o(0)
       , fabric_fpga_bid_axi_m1_o2                   =>  fabric_fpga_bid_axi_m1_o(1)
       , fabric_fpga_bid_axi_m1_o3                   =>  fabric_fpga_bid_axi_m1_o(2)
       , fabric_fpga_bid_axi_m1_o4                   =>  fabric_fpga_bid_axi_m1_o(3)
       , fabric_fpga_bid_axi_m1_o5                   =>  fabric_fpga_bid_axi_m1_o(4)
       , fabric_fpga_bresp_axi_m1_o1                 =>  fabric_fpga_bresp_axi_m1_o(0)
       , fabric_fpga_bresp_axi_m1_o2                 =>  fabric_fpga_bresp_axi_m1_o(1)
       , fabric_fpga_bvalid_axi_m1_o                 =>  fabric_fpga_bvalid_axi_m1_o
       , fabric_fpga_dma_ack_m1_o1                   =>  fabric_fpga_dma_ack_m1_o(0)
       , fabric_fpga_dma_ack_m1_o2                   =>  fabric_fpga_dma_ack_m1_o(1)
       , fabric_fpga_dma_ack_m1_o3                   =>  fabric_fpga_dma_ack_m1_o(2)
       , fabric_fpga_dma_ack_m1_o4                   =>  fabric_fpga_dma_ack_m1_o(3)
       , fabric_fpga_dma_ack_m1_o5                   =>  fabric_fpga_dma_ack_m1_o(4)
       , fabric_fpga_dma_ack_m1_o6                   =>  fabric_fpga_dma_ack_m1_o(5)
       , fabric_fpga_dma_finish_m1_o1                =>  fabric_fpga_dma_finish_m1_o(0)
       , fabric_fpga_dma_finish_m1_o2                =>  fabric_fpga_dma_finish_m1_o(1)
       , fabric_fpga_dma_finish_m1_o3                =>  fabric_fpga_dma_finish_m1_o(2)
       , fabric_fpga_dma_finish_m1_o4                =>  fabric_fpga_dma_finish_m1_o(3)
       , fabric_fpga_dma_finish_m1_o5                =>  fabric_fpga_dma_finish_m1_o(4)
       , fabric_fpga_dma_finish_m1_o6                =>  fabric_fpga_dma_finish_m1_o(5)
       , fabric_fpga_rdata_axi_m1_o1                 =>  fabric_fpga_rdata_axi_m1_o(0)
       , fabric_fpga_rdata_axi_m1_o2                 =>  fabric_fpga_rdata_axi_m1_o(1)
       , fabric_fpga_rdata_axi_m1_o3                 =>  fabric_fpga_rdata_axi_m1_o(2)
       , fabric_fpga_rdata_axi_m1_o4                 =>  fabric_fpga_rdata_axi_m1_o(3)
       , fabric_fpga_rdata_axi_m1_o5                 =>  fabric_fpga_rdata_axi_m1_o(4)
       , fabric_fpga_rdata_axi_m1_o6                 =>  fabric_fpga_rdata_axi_m1_o(5)
       , fabric_fpga_rdata_axi_m1_o7                 =>  fabric_fpga_rdata_axi_m1_o(6)
       , fabric_fpga_rdata_axi_m1_o8                 =>  fabric_fpga_rdata_axi_m1_o(7)
       , fabric_fpga_rdata_axi_m1_o9                 =>  fabric_fpga_rdata_axi_m1_o(8)
       , fabric_fpga_rdata_axi_m1_o10                =>  fabric_fpga_rdata_axi_m1_o(9)
       , fabric_fpga_rdata_axi_m1_o11                =>  fabric_fpga_rdata_axi_m1_o(10)
       , fabric_fpga_rdata_axi_m1_o12                =>  fabric_fpga_rdata_axi_m1_o(11)
       , fabric_fpga_rdata_axi_m1_o13                =>  fabric_fpga_rdata_axi_m1_o(12)
       , fabric_fpga_rdata_axi_m1_o14                =>  fabric_fpga_rdata_axi_m1_o(13)
       , fabric_fpga_rdata_axi_m1_o15                =>  fabric_fpga_rdata_axi_m1_o(14)
       , fabric_fpga_rdata_axi_m1_o16                =>  fabric_fpga_rdata_axi_m1_o(15)
       , fabric_fpga_rdata_axi_m1_o17                =>  fabric_fpga_rdata_axi_m1_o(16)
       , fabric_fpga_rdata_axi_m1_o18                =>  fabric_fpga_rdata_axi_m1_o(17)
       , fabric_fpga_rdata_axi_m1_o19                =>  fabric_fpga_rdata_axi_m1_o(18)
       , fabric_fpga_rdata_axi_m1_o20                =>  fabric_fpga_rdata_axi_m1_o(19)
       , fabric_fpga_rdata_axi_m1_o21                =>  fabric_fpga_rdata_axi_m1_o(20)
       , fabric_fpga_rdata_axi_m1_o22                =>  fabric_fpga_rdata_axi_m1_o(21)
       , fabric_fpga_rdata_axi_m1_o23                =>  fabric_fpga_rdata_axi_m1_o(22)
       , fabric_fpga_rdata_axi_m1_o24                =>  fabric_fpga_rdata_axi_m1_o(23)
       , fabric_fpga_rdata_axi_m1_o25                =>  fabric_fpga_rdata_axi_m1_o(24)
       , fabric_fpga_rdata_axi_m1_o26                =>  fabric_fpga_rdata_axi_m1_o(25)
       , fabric_fpga_rdata_axi_m1_o27                =>  fabric_fpga_rdata_axi_m1_o(26)
       , fabric_fpga_rdata_axi_m1_o28                =>  fabric_fpga_rdata_axi_m1_o(27)
       , fabric_fpga_rdata_axi_m1_o29                =>  fabric_fpga_rdata_axi_m1_o(28)
       , fabric_fpga_rdata_axi_m1_o30                =>  fabric_fpga_rdata_axi_m1_o(29)
       , fabric_fpga_rdata_axi_m1_o31                =>  fabric_fpga_rdata_axi_m1_o(30)
       , fabric_fpga_rdata_axi_m1_o32                =>  fabric_fpga_rdata_axi_m1_o(31)
       , fabric_fpga_rdata_axi_m1_o33                =>  fabric_fpga_rdata_axi_m1_o(32)
       , fabric_fpga_rdata_axi_m1_o34                =>  fabric_fpga_rdata_axi_m1_o(33)
       , fabric_fpga_rdata_axi_m1_o35                =>  fabric_fpga_rdata_axi_m1_o(34)
       , fabric_fpga_rdata_axi_m1_o36                =>  fabric_fpga_rdata_axi_m1_o(35)
       , fabric_fpga_rdata_axi_m1_o37                =>  fabric_fpga_rdata_axi_m1_o(36)
       , fabric_fpga_rdata_axi_m1_o38                =>  fabric_fpga_rdata_axi_m1_o(37)
       , fabric_fpga_rdata_axi_m1_o39                =>  fabric_fpga_rdata_axi_m1_o(38)
       , fabric_fpga_rdata_axi_m1_o40                =>  fabric_fpga_rdata_axi_m1_o(39)
       , fabric_fpga_rdata_axi_m1_o41                =>  fabric_fpga_rdata_axi_m1_o(40)
       , fabric_fpga_rdata_axi_m1_o42                =>  fabric_fpga_rdata_axi_m1_o(41)
       , fabric_fpga_rdata_axi_m1_o43                =>  fabric_fpga_rdata_axi_m1_o(42)
       , fabric_fpga_rdata_axi_m1_o44                =>  fabric_fpga_rdata_axi_m1_o(43)
       , fabric_fpga_rdata_axi_m1_o45                =>  fabric_fpga_rdata_axi_m1_o(44)
       , fabric_fpga_rdata_axi_m1_o46                =>  fabric_fpga_rdata_axi_m1_o(45)
       , fabric_fpga_rdata_axi_m1_o47                =>  fabric_fpga_rdata_axi_m1_o(46)
       , fabric_fpga_rdata_axi_m1_o48                =>  fabric_fpga_rdata_axi_m1_o(47)
       , fabric_fpga_rdata_axi_m1_o49                =>  fabric_fpga_rdata_axi_m1_o(48)
       , fabric_fpga_rdata_axi_m1_o50                =>  fabric_fpga_rdata_axi_m1_o(49)
       , fabric_fpga_rdata_axi_m1_o51                =>  fabric_fpga_rdata_axi_m1_o(50)
       , fabric_fpga_rdata_axi_m1_o52                =>  fabric_fpga_rdata_axi_m1_o(51)
       , fabric_fpga_rdata_axi_m1_o53                =>  fabric_fpga_rdata_axi_m1_o(52)
       , fabric_fpga_rdata_axi_m1_o54                =>  fabric_fpga_rdata_axi_m1_o(53)
       , fabric_fpga_rdata_axi_m1_o55                =>  fabric_fpga_rdata_axi_m1_o(54)
       , fabric_fpga_rdata_axi_m1_o56                =>  fabric_fpga_rdata_axi_m1_o(55)
       , fabric_fpga_rdata_axi_m1_o57                =>  fabric_fpga_rdata_axi_m1_o(56)
       , fabric_fpga_rdata_axi_m1_o58                =>  fabric_fpga_rdata_axi_m1_o(57)
       , fabric_fpga_rdata_axi_m1_o59                =>  fabric_fpga_rdata_axi_m1_o(58)
       , fabric_fpga_rdata_axi_m1_o60                =>  fabric_fpga_rdata_axi_m1_o(59)
       , fabric_fpga_rdata_axi_m1_o61                =>  fabric_fpga_rdata_axi_m1_o(60)
       , fabric_fpga_rdata_axi_m1_o62                =>  fabric_fpga_rdata_axi_m1_o(61)
       , fabric_fpga_rdata_axi_m1_o63                =>  fabric_fpga_rdata_axi_m1_o(62)
       , fabric_fpga_rdata_axi_m1_o64                =>  fabric_fpga_rdata_axi_m1_o(63)
       , fabric_fpga_rdata_axi_m1_o65                =>  fabric_fpga_rdata_axi_m1_o(64)
       , fabric_fpga_rdata_axi_m1_o66                =>  fabric_fpga_rdata_axi_m1_o(65)
       , fabric_fpga_rdata_axi_m1_o67                =>  fabric_fpga_rdata_axi_m1_o(66)
       , fabric_fpga_rdata_axi_m1_o68                =>  fabric_fpga_rdata_axi_m1_o(67)
       , fabric_fpga_rdata_axi_m1_o69                =>  fabric_fpga_rdata_axi_m1_o(68)
       , fabric_fpga_rdata_axi_m1_o70                =>  fabric_fpga_rdata_axi_m1_o(69)
       , fabric_fpga_rdata_axi_m1_o71                =>  fabric_fpga_rdata_axi_m1_o(70)
       , fabric_fpga_rdata_axi_m1_o72                =>  fabric_fpga_rdata_axi_m1_o(71)
       , fabric_fpga_rdata_axi_m1_o73                =>  fabric_fpga_rdata_axi_m1_o(72)
       , fabric_fpga_rdata_axi_m1_o74                =>  fabric_fpga_rdata_axi_m1_o(73)
       , fabric_fpga_rdata_axi_m1_o75                =>  fabric_fpga_rdata_axi_m1_o(74)
       , fabric_fpga_rdata_axi_m1_o76                =>  fabric_fpga_rdata_axi_m1_o(75)
       , fabric_fpga_rdata_axi_m1_o77                =>  fabric_fpga_rdata_axi_m1_o(76)
       , fabric_fpga_rdata_axi_m1_o78                =>  fabric_fpga_rdata_axi_m1_o(77)
       , fabric_fpga_rdata_axi_m1_o79                =>  fabric_fpga_rdata_axi_m1_o(78)
       , fabric_fpga_rdata_axi_m1_o80                =>  fabric_fpga_rdata_axi_m1_o(79)
       , fabric_fpga_rdata_axi_m1_o81                =>  fabric_fpga_rdata_axi_m1_o(80)
       , fabric_fpga_rdata_axi_m1_o82                =>  fabric_fpga_rdata_axi_m1_o(81)
       , fabric_fpga_rdata_axi_m1_o83                =>  fabric_fpga_rdata_axi_m1_o(82)
       , fabric_fpga_rdata_axi_m1_o84                =>  fabric_fpga_rdata_axi_m1_o(83)
       , fabric_fpga_rdata_axi_m1_o85                =>  fabric_fpga_rdata_axi_m1_o(84)
       , fabric_fpga_rdata_axi_m1_o86                =>  fabric_fpga_rdata_axi_m1_o(85)
       , fabric_fpga_rdata_axi_m1_o87                =>  fabric_fpga_rdata_axi_m1_o(86)
       , fabric_fpga_rdata_axi_m1_o88                =>  fabric_fpga_rdata_axi_m1_o(87)
       , fabric_fpga_rdata_axi_m1_o89                =>  fabric_fpga_rdata_axi_m1_o(88)
       , fabric_fpga_rdata_axi_m1_o90                =>  fabric_fpga_rdata_axi_m1_o(89)
       , fabric_fpga_rdata_axi_m1_o91                =>  fabric_fpga_rdata_axi_m1_o(90)
       , fabric_fpga_rdata_axi_m1_o92                =>  fabric_fpga_rdata_axi_m1_o(91)
       , fabric_fpga_rdata_axi_m1_o93                =>  fabric_fpga_rdata_axi_m1_o(92)
       , fabric_fpga_rdata_axi_m1_o94                =>  fabric_fpga_rdata_axi_m1_o(93)
       , fabric_fpga_rdata_axi_m1_o95                =>  fabric_fpga_rdata_axi_m1_o(94)
       , fabric_fpga_rdata_axi_m1_o96                =>  fabric_fpga_rdata_axi_m1_o(95)
       , fabric_fpga_rdata_axi_m1_o97                =>  fabric_fpga_rdata_axi_m1_o(96)
       , fabric_fpga_rdata_axi_m1_o98                =>  fabric_fpga_rdata_axi_m1_o(97)
       , fabric_fpga_rdata_axi_m1_o99                =>  fabric_fpga_rdata_axi_m1_o(98)
       , fabric_fpga_rdata_axi_m1_o100               =>  fabric_fpga_rdata_axi_m1_o(99)
       , fabric_fpga_rdata_axi_m1_o101               =>  fabric_fpga_rdata_axi_m1_o(100)
       , fabric_fpga_rdata_axi_m1_o102               =>  fabric_fpga_rdata_axi_m1_o(101)
       , fabric_fpga_rdata_axi_m1_o103               =>  fabric_fpga_rdata_axi_m1_o(102)
       , fabric_fpga_rdata_axi_m1_o104               =>  fabric_fpga_rdata_axi_m1_o(103)
       , fabric_fpga_rdata_axi_m1_o105               =>  fabric_fpga_rdata_axi_m1_o(104)
       , fabric_fpga_rdata_axi_m1_o106               =>  fabric_fpga_rdata_axi_m1_o(105)
       , fabric_fpga_rdata_axi_m1_o107               =>  fabric_fpga_rdata_axi_m1_o(106)
       , fabric_fpga_rdata_axi_m1_o108               =>  fabric_fpga_rdata_axi_m1_o(107)
       , fabric_fpga_rdata_axi_m1_o109               =>  fabric_fpga_rdata_axi_m1_o(108)
       , fabric_fpga_rdata_axi_m1_o110               =>  fabric_fpga_rdata_axi_m1_o(109)
       , fabric_fpga_rdata_axi_m1_o111               =>  fabric_fpga_rdata_axi_m1_o(110)
       , fabric_fpga_rdata_axi_m1_o112               =>  fabric_fpga_rdata_axi_m1_o(111)
       , fabric_fpga_rdata_axi_m1_o113               =>  fabric_fpga_rdata_axi_m1_o(112)
       , fabric_fpga_rdata_axi_m1_o114               =>  fabric_fpga_rdata_axi_m1_o(113)
       , fabric_fpga_rdata_axi_m1_o115               =>  fabric_fpga_rdata_axi_m1_o(114)
       , fabric_fpga_rdata_axi_m1_o116               =>  fabric_fpga_rdata_axi_m1_o(115)
       , fabric_fpga_rdata_axi_m1_o117               =>  fabric_fpga_rdata_axi_m1_o(116)
       , fabric_fpga_rdata_axi_m1_o118               =>  fabric_fpga_rdata_axi_m1_o(117)
       , fabric_fpga_rdata_axi_m1_o119               =>  fabric_fpga_rdata_axi_m1_o(118)
       , fabric_fpga_rdata_axi_m1_o120               =>  fabric_fpga_rdata_axi_m1_o(119)
       , fabric_fpga_rdata_axi_m1_o121               =>  fabric_fpga_rdata_axi_m1_o(120)
       , fabric_fpga_rdata_axi_m1_o122               =>  fabric_fpga_rdata_axi_m1_o(121)
       , fabric_fpga_rdata_axi_m1_o123               =>  fabric_fpga_rdata_axi_m1_o(122)
       , fabric_fpga_rdata_axi_m1_o124               =>  fabric_fpga_rdata_axi_m1_o(123)
       , fabric_fpga_rdata_axi_m1_o125               =>  fabric_fpga_rdata_axi_m1_o(124)
       , fabric_fpga_rdata_axi_m1_o126               =>  fabric_fpga_rdata_axi_m1_o(125)
       , fabric_fpga_rdata_axi_m1_o127               =>  fabric_fpga_rdata_axi_m1_o(126)
       , fabric_fpga_rdata_axi_m1_o128               =>  fabric_fpga_rdata_axi_m1_o(127)
       , fabric_fpga_rid_axi_m1_o1                   =>  fabric_fpga_rid_axi_m1_o(0)
       , fabric_fpga_rid_axi_m1_o2                   =>  fabric_fpga_rid_axi_m1_o(1)
       , fabric_fpga_rid_axi_m1_o3                   =>  fabric_fpga_rid_axi_m1_o(2)
       , fabric_fpga_rid_axi_m1_o4                   =>  fabric_fpga_rid_axi_m1_o(3)
       , fabric_fpga_rid_axi_m1_o5                   =>  fabric_fpga_rid_axi_m1_o(4)
       , fabric_fpga_rlast_axi_m1_o                  =>  fabric_fpga_rlast_axi_m1_o
       , fabric_fpga_rresp_axi_m1_o1                 =>  fabric_fpga_rresp_axi_m1_o(0)
       , fabric_fpga_rresp_axi_m1_o2                 =>  fabric_fpga_rresp_axi_m1_o(1)
       , fabric_fpga_rvalid_axi_m1_o                 =>  fabric_fpga_rvalid_axi_m1_o
       , fabric_fpga_wready_axi_m1_o                 =>  fabric_fpga_wready_axi_m1_o
       , fabric_fpga_araddr_axi_m1_i1                =>  fabric_fpga_araddr_axi_m1_i(0)
       , fabric_fpga_araddr_axi_m1_i2                =>  fabric_fpga_araddr_axi_m1_i(1)
       , fabric_fpga_araddr_axi_m1_i3                =>  fabric_fpga_araddr_axi_m1_i(2)
       , fabric_fpga_araddr_axi_m1_i4                =>  fabric_fpga_araddr_axi_m1_i(3)
       , fabric_fpga_araddr_axi_m1_i5                =>  fabric_fpga_araddr_axi_m1_i(4)
       , fabric_fpga_araddr_axi_m1_i6                =>  fabric_fpga_araddr_axi_m1_i(5)
       , fabric_fpga_araddr_axi_m1_i7                =>  fabric_fpga_araddr_axi_m1_i(6)
       , fabric_fpga_araddr_axi_m1_i8                =>  fabric_fpga_araddr_axi_m1_i(7)
       , fabric_fpga_araddr_axi_m1_i9                =>  fabric_fpga_araddr_axi_m1_i(8)
       , fabric_fpga_araddr_axi_m1_i10               =>  fabric_fpga_araddr_axi_m1_i(9)
       , fabric_fpga_araddr_axi_m1_i11               =>  fabric_fpga_araddr_axi_m1_i(10)
       , fabric_fpga_araddr_axi_m1_i12               =>  fabric_fpga_araddr_axi_m1_i(11)
       , fabric_fpga_araddr_axi_m1_i13               =>  fabric_fpga_araddr_axi_m1_i(12)
       , fabric_fpga_araddr_axi_m1_i14               =>  fabric_fpga_araddr_axi_m1_i(13)
       , fabric_fpga_araddr_axi_m1_i15               =>  fabric_fpga_araddr_axi_m1_i(14)
       , fabric_fpga_araddr_axi_m1_i16               =>  fabric_fpga_araddr_axi_m1_i(15)
       , fabric_fpga_araddr_axi_m1_i17               =>  fabric_fpga_araddr_axi_m1_i(16)
       , fabric_fpga_araddr_axi_m1_i18               =>  fabric_fpga_araddr_axi_m1_i(17)
       , fabric_fpga_araddr_axi_m1_i19               =>  fabric_fpga_araddr_axi_m1_i(18)
       , fabric_fpga_araddr_axi_m1_i20               =>  fabric_fpga_araddr_axi_m1_i(19)
       , fabric_fpga_araddr_axi_m1_i21               =>  fabric_fpga_araddr_axi_m1_i(20)
       , fabric_fpga_araddr_axi_m1_i22               =>  fabric_fpga_araddr_axi_m1_i(21)
       , fabric_fpga_araddr_axi_m1_i23               =>  fabric_fpga_araddr_axi_m1_i(22)
       , fabric_fpga_araddr_axi_m1_i24               =>  fabric_fpga_araddr_axi_m1_i(23)
       , fabric_fpga_araddr_axi_m1_i25               =>  fabric_fpga_araddr_axi_m1_i(24)
       , fabric_fpga_araddr_axi_m1_i26               =>  fabric_fpga_araddr_axi_m1_i(25)
       , fabric_fpga_araddr_axi_m1_i27               =>  fabric_fpga_araddr_axi_m1_i(26)
       , fabric_fpga_araddr_axi_m1_i28               =>  fabric_fpga_araddr_axi_m1_i(27)
       , fabric_fpga_araddr_axi_m1_i29               =>  fabric_fpga_araddr_axi_m1_i(28)
       , fabric_fpga_araddr_axi_m1_i30               =>  fabric_fpga_araddr_axi_m1_i(29)
       , fabric_fpga_araddr_axi_m1_i31               =>  fabric_fpga_araddr_axi_m1_i(30)
       , fabric_fpga_araddr_axi_m1_i32               =>  fabric_fpga_araddr_axi_m1_i(31)
       , fabric_fpga_araddr_axi_m1_i33               =>  fabric_fpga_araddr_axi_m1_i(32)
       , fabric_fpga_araddr_axi_m1_i34               =>  fabric_fpga_araddr_axi_m1_i(33)
       , fabric_fpga_araddr_axi_m1_i35               =>  fabric_fpga_araddr_axi_m1_i(34)
       , fabric_fpga_araddr_axi_m1_i36               =>  fabric_fpga_araddr_axi_m1_i(35)
       , fabric_fpga_araddr_axi_m1_i37               =>  fabric_fpga_araddr_axi_m1_i(36)
       , fabric_fpga_araddr_axi_m1_i38               =>  fabric_fpga_araddr_axi_m1_i(37)
       , fabric_fpga_araddr_axi_m1_i39               =>  fabric_fpga_araddr_axi_m1_i(38)
       , fabric_fpga_araddr_axi_m1_i40               =>  fabric_fpga_araddr_axi_m1_i(39)
       , fabric_fpga_arburst_axi_m1_i1               =>  fabric_fpga_arburst_axi_m1_i(0)
       , fabric_fpga_arburst_axi_m1_i2               =>  fabric_fpga_arburst_axi_m1_i(1)
       , fabric_fpga_arcache_axi_m1_i1               =>  fabric_fpga_arcache_axi_m1_i(0)
       , fabric_fpga_arcache_axi_m1_i2               =>  fabric_fpga_arcache_axi_m1_i(1)
       , fabric_fpga_arcache_axi_m1_i3               =>  fabric_fpga_arcache_axi_m1_i(2)
       , fabric_fpga_arcache_axi_m1_i4               =>  fabric_fpga_arcache_axi_m1_i(3)
       , fabric_fpga_arid_axi_m1_i1                  =>  fabric_fpga_arid_axi_m1_i(0)
       , fabric_fpga_arid_axi_m1_i2                  =>  fabric_fpga_arid_axi_m1_i(1)
       , fabric_fpga_arid_axi_m1_i3                  =>  fabric_fpga_arid_axi_m1_i(2)
       , fabric_fpga_arid_axi_m1_i4                  =>  fabric_fpga_arid_axi_m1_i(3)
       , fabric_fpga_arid_axi_m1_i5                  =>  fabric_fpga_arid_axi_m1_i(4)
       , fabric_fpga_arlen_axi_m1_i1                 =>  fabric_fpga_arlen_axi_m1_i(0)
       , fabric_fpga_arlen_axi_m1_i2                 =>  fabric_fpga_arlen_axi_m1_i(1)
       , fabric_fpga_arlen_axi_m1_i3                 =>  fabric_fpga_arlen_axi_m1_i(2)
       , fabric_fpga_arlen_axi_m1_i4                 =>  fabric_fpga_arlen_axi_m1_i(3)
       , fabric_fpga_arlen_axi_m1_i5                 =>  fabric_fpga_arlen_axi_m1_i(4)
       , fabric_fpga_arlen_axi_m1_i6                 =>  fabric_fpga_arlen_axi_m1_i(5)
       , fabric_fpga_arlen_axi_m1_i7                 =>  fabric_fpga_arlen_axi_m1_i(6)
       , fabric_fpga_arlen_axi_m1_i8                 =>  fabric_fpga_arlen_axi_m1_i(7)
       , fabric_fpga_arlock_axi_m1_i                 =>  fabric_fpga_arlock_axi_m1_i
       , fabric_fpga_arprot_axi_m1_i1                =>  fabric_fpga_arprot_axi_m1_i(0)
       , fabric_fpga_arprot_axi_m1_i2                =>  fabric_fpga_arprot_axi_m1_i(1)
       , fabric_fpga_arprot_axi_m1_i3                =>  fabric_fpga_arprot_axi_m1_i(2)
       , fabric_fpga_arqos_axi_m1_i1                 =>  fabric_fpga_arqos_axi_m1_i(0)
       , fabric_fpga_arqos_axi_m1_i2                 =>  fabric_fpga_arqos_axi_m1_i(1)
       , fabric_fpga_arqos_axi_m1_i3                 =>  fabric_fpga_arqos_axi_m1_i(2)
       , fabric_fpga_arqos_axi_m1_i4                 =>  fabric_fpga_arqos_axi_m1_i(3)
       , fabric_fpga_arsize_axi_m1_i1                =>  fabric_fpga_arsize_axi_m1_i(0)
       , fabric_fpga_arsize_axi_m1_i2                =>  fabric_fpga_arsize_axi_m1_i(1)
       , fabric_fpga_arsize_axi_m1_i3                =>  fabric_fpga_arsize_axi_m1_i(2)
       , fabric_fpga_arvalid_axi_m1_i                =>  fabric_fpga_arvalid_axi_m1_i
       , fabric_fpga_awaddr_axi_m1_i1                =>  fabric_fpga_awaddr_axi_m1_i(0)
       , fabric_fpga_awaddr_axi_m1_i2                =>  fabric_fpga_awaddr_axi_m1_i(1)
       , fabric_fpga_awaddr_axi_m1_i3                =>  fabric_fpga_awaddr_axi_m1_i(2)
       , fabric_fpga_awaddr_axi_m1_i4                =>  fabric_fpga_awaddr_axi_m1_i(3)
       , fabric_fpga_awaddr_axi_m1_i5                =>  fabric_fpga_awaddr_axi_m1_i(4)
       , fabric_fpga_awaddr_axi_m1_i6                =>  fabric_fpga_awaddr_axi_m1_i(5)
       , fabric_fpga_awaddr_axi_m1_i7                =>  fabric_fpga_awaddr_axi_m1_i(6)
       , fabric_fpga_awaddr_axi_m1_i8                =>  fabric_fpga_awaddr_axi_m1_i(7)
       , fabric_fpga_awaddr_axi_m1_i9                =>  fabric_fpga_awaddr_axi_m1_i(8)
       , fabric_fpga_awaddr_axi_m1_i10               =>  fabric_fpga_awaddr_axi_m1_i(9)
       , fabric_fpga_awaddr_axi_m1_i11               =>  fabric_fpga_awaddr_axi_m1_i(10)
       , fabric_fpga_awaddr_axi_m1_i12               =>  fabric_fpga_awaddr_axi_m1_i(11)
       , fabric_fpga_awaddr_axi_m1_i13               =>  fabric_fpga_awaddr_axi_m1_i(12)
       , fabric_fpga_awaddr_axi_m1_i14               =>  fabric_fpga_awaddr_axi_m1_i(13)
       , fabric_fpga_awaddr_axi_m1_i15               =>  fabric_fpga_awaddr_axi_m1_i(14)
       , fabric_fpga_awaddr_axi_m1_i16               =>  fabric_fpga_awaddr_axi_m1_i(15)
       , fabric_fpga_awaddr_axi_m1_i17               =>  fabric_fpga_awaddr_axi_m1_i(16)
       , fabric_fpga_awaddr_axi_m1_i18               =>  fabric_fpga_awaddr_axi_m1_i(17)
       , fabric_fpga_awaddr_axi_m1_i19               =>  fabric_fpga_awaddr_axi_m1_i(18)
       , fabric_fpga_awaddr_axi_m1_i20               =>  fabric_fpga_awaddr_axi_m1_i(19)
       , fabric_fpga_awaddr_axi_m1_i21               =>  fabric_fpga_awaddr_axi_m1_i(20)
       , fabric_fpga_awaddr_axi_m1_i22               =>  fabric_fpga_awaddr_axi_m1_i(21)
       , fabric_fpga_awaddr_axi_m1_i23               =>  fabric_fpga_awaddr_axi_m1_i(22)
       , fabric_fpga_awaddr_axi_m1_i24               =>  fabric_fpga_awaddr_axi_m1_i(23)
       , fabric_fpga_awaddr_axi_m1_i25               =>  fabric_fpga_awaddr_axi_m1_i(24)
       , fabric_fpga_awaddr_axi_m1_i26               =>  fabric_fpga_awaddr_axi_m1_i(25)
       , fabric_fpga_awaddr_axi_m1_i27               =>  fabric_fpga_awaddr_axi_m1_i(26)
       , fabric_fpga_awaddr_axi_m1_i28               =>  fabric_fpga_awaddr_axi_m1_i(27)
       , fabric_fpga_awaddr_axi_m1_i29               =>  fabric_fpga_awaddr_axi_m1_i(28)
       , fabric_fpga_awaddr_axi_m1_i30               =>  fabric_fpga_awaddr_axi_m1_i(29)
       , fabric_fpga_awaddr_axi_m1_i31               =>  fabric_fpga_awaddr_axi_m1_i(30)
       , fabric_fpga_awaddr_axi_m1_i32               =>  fabric_fpga_awaddr_axi_m1_i(31)
       , fabric_fpga_awaddr_axi_m1_i33               =>  fabric_fpga_awaddr_axi_m1_i(32)
       , fabric_fpga_awaddr_axi_m1_i34               =>  fabric_fpga_awaddr_axi_m1_i(33)
       , fabric_fpga_awaddr_axi_m1_i35               =>  fabric_fpga_awaddr_axi_m1_i(34)
       , fabric_fpga_awaddr_axi_m1_i36               =>  fabric_fpga_awaddr_axi_m1_i(35)
       , fabric_fpga_awaddr_axi_m1_i37               =>  fabric_fpga_awaddr_axi_m1_i(36)
       , fabric_fpga_awaddr_axi_m1_i38               =>  fabric_fpga_awaddr_axi_m1_i(37)
       , fabric_fpga_awaddr_axi_m1_i39               =>  fabric_fpga_awaddr_axi_m1_i(38)
       , fabric_fpga_awaddr_axi_m1_i40               =>  fabric_fpga_awaddr_axi_m1_i(39)
       , fabric_fpga_awburst_axi_m1_i1               =>  fabric_fpga_awburst_axi_m1_i(0)
       , fabric_fpga_awburst_axi_m1_i2               =>  fabric_fpga_awburst_axi_m1_i(1)
       , fabric_fpga_awcache_axi_m1_i1               =>  fabric_fpga_awcache_axi_m1_i(0)
       , fabric_fpga_awcache_axi_m1_i2               =>  fabric_fpga_awcache_axi_m1_i(1)
       , fabric_fpga_awcache_axi_m1_i3               =>  fabric_fpga_awcache_axi_m1_i(2)
       , fabric_fpga_awcache_axi_m1_i4               =>  fabric_fpga_awcache_axi_m1_i(3)
       , fabric_fpga_awid_axi_m1_i1                  =>  fabric_fpga_awid_axi_m1_i(0)
       , fabric_fpga_awid_axi_m1_i2                  =>  fabric_fpga_awid_axi_m1_i(1)
       , fabric_fpga_awid_axi_m1_i3                  =>  fabric_fpga_awid_axi_m1_i(2)
       , fabric_fpga_awid_axi_m1_i4                  =>  fabric_fpga_awid_axi_m1_i(3)
       , fabric_fpga_awid_axi_m1_i5                  =>  fabric_fpga_awid_axi_m1_i(4)
       , fabric_fpga_awlen_axi_m1_i1                 =>  fabric_fpga_awlen_axi_m1_i(0)
       , fabric_fpga_awlen_axi_m1_i2                 =>  fabric_fpga_awlen_axi_m1_i(1)
       , fabric_fpga_awlen_axi_m1_i3                 =>  fabric_fpga_awlen_axi_m1_i(2)
       , fabric_fpga_awlen_axi_m1_i4                 =>  fabric_fpga_awlen_axi_m1_i(3)
       , fabric_fpga_awlen_axi_m1_i5                 =>  fabric_fpga_awlen_axi_m1_i(4)
       , fabric_fpga_awlen_axi_m1_i6                 =>  fabric_fpga_awlen_axi_m1_i(5)
       , fabric_fpga_awlen_axi_m1_i7                 =>  fabric_fpga_awlen_axi_m1_i(6)
       , fabric_fpga_awlen_axi_m1_i8                 =>  fabric_fpga_awlen_axi_m1_i(7)
       , fabric_fpga_awlock_axi_m1_i                 =>  fabric_fpga_awlock_axi_m1_i
       , fabric_fpga_awprot_axi_m1_i1                =>  fabric_fpga_awprot_axi_m1_i(0)
       , fabric_fpga_awprot_axi_m1_i2                =>  fabric_fpga_awprot_axi_m1_i(1)
       , fabric_fpga_awprot_axi_m1_i3                =>  fabric_fpga_awprot_axi_m1_i(2)
       , fabric_fpga_awqos_axi_m1_i1                 =>  fabric_fpga_awqos_axi_m1_i(0)
       , fabric_fpga_awqos_axi_m1_i2                 =>  fabric_fpga_awqos_axi_m1_i(1)
       , fabric_fpga_awqos_axi_m1_i3                 =>  fabric_fpga_awqos_axi_m1_i(2)
       , fabric_fpga_awqos_axi_m1_i4                 =>  fabric_fpga_awqos_axi_m1_i(3)
       , fabric_fpga_awsize_axi_m1_i1                =>  fabric_fpga_awsize_axi_m1_i(0)
       , fabric_fpga_awsize_axi_m1_i2                =>  fabric_fpga_awsize_axi_m1_i(1)
       , fabric_fpga_awsize_axi_m1_i3                =>  fabric_fpga_awsize_axi_m1_i(2)
       , fabric_fpga_awvalid_axi_m1_i                =>  fabric_fpga_awvalid_axi_m1_i
       , fabric_fpga_bready_axi_m1_i                 =>  fabric_fpga_bready_axi_m1_i
       , fabric_fpga_dma_last_m1_i1                  =>  fabric_fpga_dma_last_m1_i(0)
       , fabric_fpga_dma_last_m1_i2                  =>  fabric_fpga_dma_last_m1_i(1)
       , fabric_fpga_dma_last_m1_i3                  =>  fabric_fpga_dma_last_m1_i(2)
       , fabric_fpga_dma_last_m1_i4                  =>  fabric_fpga_dma_last_m1_i(3)
       , fabric_fpga_dma_last_m1_i5                  =>  fabric_fpga_dma_last_m1_i(4)
       , fabric_fpga_dma_last_m1_i6                  =>  fabric_fpga_dma_last_m1_i(5)
       , fabric_fpga_dma_req_m1_i1                   =>  fabric_fpga_dma_req_m1_i(0)
       , fabric_fpga_dma_req_m1_i2                   =>  fabric_fpga_dma_req_m1_i(1)
       , fabric_fpga_dma_req_m1_i3                   =>  fabric_fpga_dma_req_m1_i(2)
       , fabric_fpga_dma_req_m1_i4                   =>  fabric_fpga_dma_req_m1_i(3)
       , fabric_fpga_dma_req_m1_i5                   =>  fabric_fpga_dma_req_m1_i(4)
       , fabric_fpga_dma_req_m1_i6                   =>  fabric_fpga_dma_req_m1_i(5)
       , fabric_fpga_dma_single_m1_i1                =>  fabric_fpga_dma_single_m1_i(0)
       , fabric_fpga_dma_single_m1_i2                =>  fabric_fpga_dma_single_m1_i(1)
       , fabric_fpga_dma_single_m1_i3                =>  fabric_fpga_dma_single_m1_i(2)
       , fabric_fpga_dma_single_m1_i4                =>  fabric_fpga_dma_single_m1_i(3)
       , fabric_fpga_dma_single_m1_i5                =>  fabric_fpga_dma_single_m1_i(4)
       , fabric_fpga_dma_single_m1_i6                =>  fabric_fpga_dma_single_m1_i(5)
       , fabric_fpga_rready_axi_m1_i                 =>  fabric_fpga_rready_axi_m1_i
       , fabric_fpga_wdata_axi_m1_i1                 =>  fabric_fpga_wdata_axi_m1_i(0)
       , fabric_fpga_wdata_axi_m1_i2                 =>  fabric_fpga_wdata_axi_m1_i(1)
       , fabric_fpga_wdata_axi_m1_i3                 =>  fabric_fpga_wdata_axi_m1_i(2)
       , fabric_fpga_wdata_axi_m1_i4                 =>  fabric_fpga_wdata_axi_m1_i(3)
       , fabric_fpga_wdata_axi_m1_i5                 =>  fabric_fpga_wdata_axi_m1_i(4)
       , fabric_fpga_wdata_axi_m1_i6                 =>  fabric_fpga_wdata_axi_m1_i(5)
       , fabric_fpga_wdata_axi_m1_i7                 =>  fabric_fpga_wdata_axi_m1_i(6)
       , fabric_fpga_wdata_axi_m1_i8                 =>  fabric_fpga_wdata_axi_m1_i(7)
       , fabric_fpga_wdata_axi_m1_i9                 =>  fabric_fpga_wdata_axi_m1_i(8)
       , fabric_fpga_wdata_axi_m1_i10                =>  fabric_fpga_wdata_axi_m1_i(9)
       , fabric_fpga_wdata_axi_m1_i11                =>  fabric_fpga_wdata_axi_m1_i(10)
       , fabric_fpga_wdata_axi_m1_i12                =>  fabric_fpga_wdata_axi_m1_i(11)
       , fabric_fpga_wdata_axi_m1_i13                =>  fabric_fpga_wdata_axi_m1_i(12)
       , fabric_fpga_wdata_axi_m1_i14                =>  fabric_fpga_wdata_axi_m1_i(13)
       , fabric_fpga_wdata_axi_m1_i15                =>  fabric_fpga_wdata_axi_m1_i(14)
       , fabric_fpga_wdata_axi_m1_i16                =>  fabric_fpga_wdata_axi_m1_i(15)
       , fabric_fpga_wdata_axi_m1_i17                =>  fabric_fpga_wdata_axi_m1_i(16)
       , fabric_fpga_wdata_axi_m1_i18                =>  fabric_fpga_wdata_axi_m1_i(17)
       , fabric_fpga_wdata_axi_m1_i19                =>  fabric_fpga_wdata_axi_m1_i(18)
       , fabric_fpga_wdata_axi_m1_i20                =>  fabric_fpga_wdata_axi_m1_i(19)
       , fabric_fpga_wdata_axi_m1_i21                =>  fabric_fpga_wdata_axi_m1_i(20)
       , fabric_fpga_wdata_axi_m1_i22                =>  fabric_fpga_wdata_axi_m1_i(21)
       , fabric_fpga_wdata_axi_m1_i23                =>  fabric_fpga_wdata_axi_m1_i(22)
       , fabric_fpga_wdata_axi_m1_i24                =>  fabric_fpga_wdata_axi_m1_i(23)
       , fabric_fpga_wdata_axi_m1_i25                =>  fabric_fpga_wdata_axi_m1_i(24)
       , fabric_fpga_wdata_axi_m1_i26                =>  fabric_fpga_wdata_axi_m1_i(25)
       , fabric_fpga_wdata_axi_m1_i27                =>  fabric_fpga_wdata_axi_m1_i(26)
       , fabric_fpga_wdata_axi_m1_i28                =>  fabric_fpga_wdata_axi_m1_i(27)
       , fabric_fpga_wdata_axi_m1_i29                =>  fabric_fpga_wdata_axi_m1_i(28)
       , fabric_fpga_wdata_axi_m1_i30                =>  fabric_fpga_wdata_axi_m1_i(29)
       , fabric_fpga_wdata_axi_m1_i31                =>  fabric_fpga_wdata_axi_m1_i(30)
       , fabric_fpga_wdata_axi_m1_i32                =>  fabric_fpga_wdata_axi_m1_i(31)
       , fabric_fpga_wdata_axi_m1_i33                =>  fabric_fpga_wdata_axi_m1_i(32)
       , fabric_fpga_wdata_axi_m1_i34                =>  fabric_fpga_wdata_axi_m1_i(33)
       , fabric_fpga_wdata_axi_m1_i35                =>  fabric_fpga_wdata_axi_m1_i(34)
       , fabric_fpga_wdata_axi_m1_i36                =>  fabric_fpga_wdata_axi_m1_i(35)
       , fabric_fpga_wdata_axi_m1_i37                =>  fabric_fpga_wdata_axi_m1_i(36)
       , fabric_fpga_wdata_axi_m1_i38                =>  fabric_fpga_wdata_axi_m1_i(37)
       , fabric_fpga_wdata_axi_m1_i39                =>  fabric_fpga_wdata_axi_m1_i(38)
       , fabric_fpga_wdata_axi_m1_i40                =>  fabric_fpga_wdata_axi_m1_i(39)
       , fabric_fpga_wdata_axi_m1_i41                =>  fabric_fpga_wdata_axi_m1_i(40)
       , fabric_fpga_wdata_axi_m1_i42                =>  fabric_fpga_wdata_axi_m1_i(41)
       , fabric_fpga_wdata_axi_m1_i43                =>  fabric_fpga_wdata_axi_m1_i(42)
       , fabric_fpga_wdata_axi_m1_i44                =>  fabric_fpga_wdata_axi_m1_i(43)
       , fabric_fpga_wdata_axi_m1_i45                =>  fabric_fpga_wdata_axi_m1_i(44)
       , fabric_fpga_wdata_axi_m1_i46                =>  fabric_fpga_wdata_axi_m1_i(45)
       , fabric_fpga_wdata_axi_m1_i47                =>  fabric_fpga_wdata_axi_m1_i(46)
       , fabric_fpga_wdata_axi_m1_i48                =>  fabric_fpga_wdata_axi_m1_i(47)
       , fabric_fpga_wdata_axi_m1_i49                =>  fabric_fpga_wdata_axi_m1_i(48)
       , fabric_fpga_wdata_axi_m1_i50                =>  fabric_fpga_wdata_axi_m1_i(49)
       , fabric_fpga_wdata_axi_m1_i51                =>  fabric_fpga_wdata_axi_m1_i(50)
       , fabric_fpga_wdata_axi_m1_i52                =>  fabric_fpga_wdata_axi_m1_i(51)
       , fabric_fpga_wdata_axi_m1_i53                =>  fabric_fpga_wdata_axi_m1_i(52)
       , fabric_fpga_wdata_axi_m1_i54                =>  fabric_fpga_wdata_axi_m1_i(53)
       , fabric_fpga_wdata_axi_m1_i55                =>  fabric_fpga_wdata_axi_m1_i(54)
       , fabric_fpga_wdata_axi_m1_i56                =>  fabric_fpga_wdata_axi_m1_i(55)
       , fabric_fpga_wdata_axi_m1_i57                =>  fabric_fpga_wdata_axi_m1_i(56)
       , fabric_fpga_wdata_axi_m1_i58                =>  fabric_fpga_wdata_axi_m1_i(57)
       , fabric_fpga_wdata_axi_m1_i59                =>  fabric_fpga_wdata_axi_m1_i(58)
       , fabric_fpga_wdata_axi_m1_i60                =>  fabric_fpga_wdata_axi_m1_i(59)
       , fabric_fpga_wdata_axi_m1_i61                =>  fabric_fpga_wdata_axi_m1_i(60)
       , fabric_fpga_wdata_axi_m1_i62                =>  fabric_fpga_wdata_axi_m1_i(61)
       , fabric_fpga_wdata_axi_m1_i63                =>  fabric_fpga_wdata_axi_m1_i(62)
       , fabric_fpga_wdata_axi_m1_i64                =>  fabric_fpga_wdata_axi_m1_i(63)
       , fabric_fpga_wdata_axi_m1_i65                =>  fabric_fpga_wdata_axi_m1_i(64)
       , fabric_fpga_wdata_axi_m1_i66                =>  fabric_fpga_wdata_axi_m1_i(65)
       , fabric_fpga_wdata_axi_m1_i67                =>  fabric_fpga_wdata_axi_m1_i(66)
       , fabric_fpga_wdata_axi_m1_i68                =>  fabric_fpga_wdata_axi_m1_i(67)
       , fabric_fpga_wdata_axi_m1_i69                =>  fabric_fpga_wdata_axi_m1_i(68)
       , fabric_fpga_wdata_axi_m1_i70                =>  fabric_fpga_wdata_axi_m1_i(69)
       , fabric_fpga_wdata_axi_m1_i71                =>  fabric_fpga_wdata_axi_m1_i(70)
       , fabric_fpga_wdata_axi_m1_i72                =>  fabric_fpga_wdata_axi_m1_i(71)
       , fabric_fpga_wdata_axi_m1_i73                =>  fabric_fpga_wdata_axi_m1_i(72)
       , fabric_fpga_wdata_axi_m1_i74                =>  fabric_fpga_wdata_axi_m1_i(73)
       , fabric_fpga_wdata_axi_m1_i75                =>  fabric_fpga_wdata_axi_m1_i(74)
       , fabric_fpga_wdata_axi_m1_i76                =>  fabric_fpga_wdata_axi_m1_i(75)
       , fabric_fpga_wdata_axi_m1_i77                =>  fabric_fpga_wdata_axi_m1_i(76)
       , fabric_fpga_wdata_axi_m1_i78                =>  fabric_fpga_wdata_axi_m1_i(77)
       , fabric_fpga_wdata_axi_m1_i79                =>  fabric_fpga_wdata_axi_m1_i(78)
       , fabric_fpga_wdata_axi_m1_i80                =>  fabric_fpga_wdata_axi_m1_i(79)
       , fabric_fpga_wdata_axi_m1_i81                =>  fabric_fpga_wdata_axi_m1_i(80)
       , fabric_fpga_wdata_axi_m1_i82                =>  fabric_fpga_wdata_axi_m1_i(81)
       , fabric_fpga_wdata_axi_m1_i83                =>  fabric_fpga_wdata_axi_m1_i(82)
       , fabric_fpga_wdata_axi_m1_i84                =>  fabric_fpga_wdata_axi_m1_i(83)
       , fabric_fpga_wdata_axi_m1_i85                =>  fabric_fpga_wdata_axi_m1_i(84)
       , fabric_fpga_wdata_axi_m1_i86                =>  fabric_fpga_wdata_axi_m1_i(85)
       , fabric_fpga_wdata_axi_m1_i87                =>  fabric_fpga_wdata_axi_m1_i(86)
       , fabric_fpga_wdata_axi_m1_i88                =>  fabric_fpga_wdata_axi_m1_i(87)
       , fabric_fpga_wdata_axi_m1_i89                =>  fabric_fpga_wdata_axi_m1_i(88)
       , fabric_fpga_wdata_axi_m1_i90                =>  fabric_fpga_wdata_axi_m1_i(89)
       , fabric_fpga_wdata_axi_m1_i91                =>  fabric_fpga_wdata_axi_m1_i(90)
       , fabric_fpga_wdata_axi_m1_i92                =>  fabric_fpga_wdata_axi_m1_i(91)
       , fabric_fpga_wdata_axi_m1_i93                =>  fabric_fpga_wdata_axi_m1_i(92)
       , fabric_fpga_wdata_axi_m1_i94                =>  fabric_fpga_wdata_axi_m1_i(93)
       , fabric_fpga_wdata_axi_m1_i95                =>  fabric_fpga_wdata_axi_m1_i(94)
       , fabric_fpga_wdata_axi_m1_i96                =>  fabric_fpga_wdata_axi_m1_i(95)
       , fabric_fpga_wdata_axi_m1_i97                =>  fabric_fpga_wdata_axi_m1_i(96)
       , fabric_fpga_wdata_axi_m1_i98                =>  fabric_fpga_wdata_axi_m1_i(97)
       , fabric_fpga_wdata_axi_m1_i99                =>  fabric_fpga_wdata_axi_m1_i(98)
       , fabric_fpga_wdata_axi_m1_i100               =>  fabric_fpga_wdata_axi_m1_i(99)
       , fabric_fpga_wdata_axi_m1_i101               =>  fabric_fpga_wdata_axi_m1_i(100)
       , fabric_fpga_wdata_axi_m1_i102               =>  fabric_fpga_wdata_axi_m1_i(101)
       , fabric_fpga_wdata_axi_m1_i103               =>  fabric_fpga_wdata_axi_m1_i(102)
       , fabric_fpga_wdata_axi_m1_i104               =>  fabric_fpga_wdata_axi_m1_i(103)
       , fabric_fpga_wdata_axi_m1_i105               =>  fabric_fpga_wdata_axi_m1_i(104)
       , fabric_fpga_wdata_axi_m1_i106               =>  fabric_fpga_wdata_axi_m1_i(105)
       , fabric_fpga_wdata_axi_m1_i107               =>  fabric_fpga_wdata_axi_m1_i(106)
       , fabric_fpga_wdata_axi_m1_i108               =>  fabric_fpga_wdata_axi_m1_i(107)
       , fabric_fpga_wdata_axi_m1_i109               =>  fabric_fpga_wdata_axi_m1_i(108)
       , fabric_fpga_wdata_axi_m1_i110               =>  fabric_fpga_wdata_axi_m1_i(109)
       , fabric_fpga_wdata_axi_m1_i111               =>  fabric_fpga_wdata_axi_m1_i(110)
       , fabric_fpga_wdata_axi_m1_i112               =>  fabric_fpga_wdata_axi_m1_i(111)
       , fabric_fpga_wdata_axi_m1_i113               =>  fabric_fpga_wdata_axi_m1_i(112)
       , fabric_fpga_wdata_axi_m1_i114               =>  fabric_fpga_wdata_axi_m1_i(113)
       , fabric_fpga_wdata_axi_m1_i115               =>  fabric_fpga_wdata_axi_m1_i(114)
       , fabric_fpga_wdata_axi_m1_i116               =>  fabric_fpga_wdata_axi_m1_i(115)
       , fabric_fpga_wdata_axi_m1_i117               =>  fabric_fpga_wdata_axi_m1_i(116)
       , fabric_fpga_wdata_axi_m1_i118               =>  fabric_fpga_wdata_axi_m1_i(117)
       , fabric_fpga_wdata_axi_m1_i119               =>  fabric_fpga_wdata_axi_m1_i(118)
       , fabric_fpga_wdata_axi_m1_i120               =>  fabric_fpga_wdata_axi_m1_i(119)
       , fabric_fpga_wdata_axi_m1_i121               =>  fabric_fpga_wdata_axi_m1_i(120)
       , fabric_fpga_wdata_axi_m1_i122               =>  fabric_fpga_wdata_axi_m1_i(121)
       , fabric_fpga_wdata_axi_m1_i123               =>  fabric_fpga_wdata_axi_m1_i(122)
       , fabric_fpga_wdata_axi_m1_i124               =>  fabric_fpga_wdata_axi_m1_i(123)
       , fabric_fpga_wdata_axi_m1_i125               =>  fabric_fpga_wdata_axi_m1_i(124)
       , fabric_fpga_wdata_axi_m1_i126               =>  fabric_fpga_wdata_axi_m1_i(125)
       , fabric_fpga_wdata_axi_m1_i127               =>  fabric_fpga_wdata_axi_m1_i(126)
       , fabric_fpga_wdata_axi_m1_i128               =>  fabric_fpga_wdata_axi_m1_i(127)
       , fabric_fpga_wlast_axi_m1_i                  =>  fabric_fpga_wlast_axi_m1_i
       , fabric_fpga_wstrb_axi_m1_i1                 =>  fabric_fpga_wstrb_axi_m1_i(0)
       , fabric_fpga_wstrb_axi_m1_i2                 =>  fabric_fpga_wstrb_axi_m1_i(1)
       , fabric_fpga_wstrb_axi_m1_i3                 =>  fabric_fpga_wstrb_axi_m1_i(2)
       , fabric_fpga_wstrb_axi_m1_i4                 =>  fabric_fpga_wstrb_axi_m1_i(3)
       , fabric_fpga_wstrb_axi_m1_i5                 =>  fabric_fpga_wstrb_axi_m1_i(4)
       , fabric_fpga_wstrb_axi_m1_i6                 =>  fabric_fpga_wstrb_axi_m1_i(5)
       , fabric_fpga_wstrb_axi_m1_i7                 =>  fabric_fpga_wstrb_axi_m1_i(6)
       , fabric_fpga_wstrb_axi_m1_i8                 =>  fabric_fpga_wstrb_axi_m1_i(7)
       , fabric_fpga_wstrb_axi_m1_i9                 =>  fabric_fpga_wstrb_axi_m1_i(8)
       , fabric_fpga_wstrb_axi_m1_i10                =>  fabric_fpga_wstrb_axi_m1_i(9)
       , fabric_fpga_wstrb_axi_m1_i11                =>  fabric_fpga_wstrb_axi_m1_i(10)
       , fabric_fpga_wstrb_axi_m1_i12                =>  fabric_fpga_wstrb_axi_m1_i(11)
       , fabric_fpga_wstrb_axi_m1_i13                =>  fabric_fpga_wstrb_axi_m1_i(12)
       , fabric_fpga_wstrb_axi_m1_i14                =>  fabric_fpga_wstrb_axi_m1_i(13)
       , fabric_fpga_wstrb_axi_m1_i15                =>  fabric_fpga_wstrb_axi_m1_i(14)
       , fabric_fpga_wstrb_axi_m1_i16                =>  fabric_fpga_wstrb_axi_m1_i(15)
       , fabric_fpga_wvalid_axi_m1_i                 =>  fabric_fpga_wvalid_axi_m1_i
       , fabric_fpga_arready_axi_m2_o                =>  fabric_fpga_arready_axi_m2_o
       , fabric_fpga_awready_axi_m2_o                =>  fabric_fpga_awready_axi_m2_o
       , fabric_fpga_bid_axi_m2_o1                   =>  fabric_fpga_bid_axi_m2_o(0)
       , fabric_fpga_bid_axi_m2_o2                   =>  fabric_fpga_bid_axi_m2_o(1)
       , fabric_fpga_bid_axi_m2_o3                   =>  fabric_fpga_bid_axi_m2_o(2)
       , fabric_fpga_bid_axi_m2_o4                   =>  fabric_fpga_bid_axi_m2_o(3)
       , fabric_fpga_bid_axi_m2_o5                   =>  fabric_fpga_bid_axi_m2_o(4)
       , fabric_fpga_bresp_axi_m2_o1                 =>  fabric_fpga_bresp_axi_m2_o(0)
       , fabric_fpga_bresp_axi_m2_o2                 =>  fabric_fpga_bresp_axi_m2_o(1)
       , fabric_fpga_bvalid_axi_m2_o                 =>  fabric_fpga_bvalid_axi_m2_o
       , fabric_fpga_dma_ack_m2_o1                   =>  fabric_fpga_dma_ack_m2_o(0)
       , fabric_fpga_dma_ack_m2_o2                   =>  fabric_fpga_dma_ack_m2_o(1)
       , fabric_fpga_dma_ack_m2_o3                   =>  fabric_fpga_dma_ack_m2_o(2)
       , fabric_fpga_dma_ack_m2_o4                   =>  fabric_fpga_dma_ack_m2_o(3)
       , fabric_fpga_dma_ack_m2_o5                   =>  fabric_fpga_dma_ack_m2_o(4)
       , fabric_fpga_dma_ack_m2_o6                   =>  fabric_fpga_dma_ack_m2_o(5)
       , fabric_fpga_dma_finish_m2_o1                =>  fabric_fpga_dma_finish_m2_o(0)
       , fabric_fpga_dma_finish_m2_o2                =>  fabric_fpga_dma_finish_m2_o(1)
       , fabric_fpga_dma_finish_m2_o3                =>  fabric_fpga_dma_finish_m2_o(2)
       , fabric_fpga_dma_finish_m2_o4                =>  fabric_fpga_dma_finish_m2_o(3)
       , fabric_fpga_dma_finish_m2_o5                =>  fabric_fpga_dma_finish_m2_o(4)
       , fabric_fpga_dma_finish_m2_o6                =>  fabric_fpga_dma_finish_m2_o(5)
       , fabric_fpga_rdata_axi_m2_o1                 =>  fabric_fpga_rdata_axi_m2_o(0)
       , fabric_fpga_rdata_axi_m2_o2                 =>  fabric_fpga_rdata_axi_m2_o(1)
       , fabric_fpga_rdata_axi_m2_o3                 =>  fabric_fpga_rdata_axi_m2_o(2)
       , fabric_fpga_rdata_axi_m2_o4                 =>  fabric_fpga_rdata_axi_m2_o(3)
       , fabric_fpga_rdata_axi_m2_o5                 =>  fabric_fpga_rdata_axi_m2_o(4)
       , fabric_fpga_rdata_axi_m2_o6                 =>  fabric_fpga_rdata_axi_m2_o(5)
       , fabric_fpga_rdata_axi_m2_o7                 =>  fabric_fpga_rdata_axi_m2_o(6)
       , fabric_fpga_rdata_axi_m2_o8                 =>  fabric_fpga_rdata_axi_m2_o(7)
       , fabric_fpga_rdata_axi_m2_o9                 =>  fabric_fpga_rdata_axi_m2_o(8)
       , fabric_fpga_rdata_axi_m2_o10                =>  fabric_fpga_rdata_axi_m2_o(9)
       , fabric_fpga_rdata_axi_m2_o11                =>  fabric_fpga_rdata_axi_m2_o(10)
       , fabric_fpga_rdata_axi_m2_o12                =>  fabric_fpga_rdata_axi_m2_o(11)
       , fabric_fpga_rdata_axi_m2_o13                =>  fabric_fpga_rdata_axi_m2_o(12)
       , fabric_fpga_rdata_axi_m2_o14                =>  fabric_fpga_rdata_axi_m2_o(13)
       , fabric_fpga_rdata_axi_m2_o15                =>  fabric_fpga_rdata_axi_m2_o(14)
       , fabric_fpga_rdata_axi_m2_o16                =>  fabric_fpga_rdata_axi_m2_o(15)
       , fabric_fpga_rdata_axi_m2_o17                =>  fabric_fpga_rdata_axi_m2_o(16)
       , fabric_fpga_rdata_axi_m2_o18                =>  fabric_fpga_rdata_axi_m2_o(17)
       , fabric_fpga_rdata_axi_m2_o19                =>  fabric_fpga_rdata_axi_m2_o(18)
       , fabric_fpga_rdata_axi_m2_o20                =>  fabric_fpga_rdata_axi_m2_o(19)
       , fabric_fpga_rdata_axi_m2_o21                =>  fabric_fpga_rdata_axi_m2_o(20)
       , fabric_fpga_rdata_axi_m2_o22                =>  fabric_fpga_rdata_axi_m2_o(21)
       , fabric_fpga_rdata_axi_m2_o23                =>  fabric_fpga_rdata_axi_m2_o(22)
       , fabric_fpga_rdata_axi_m2_o24                =>  fabric_fpga_rdata_axi_m2_o(23)
       , fabric_fpga_rdata_axi_m2_o25                =>  fabric_fpga_rdata_axi_m2_o(24)
       , fabric_fpga_rdata_axi_m2_o26                =>  fabric_fpga_rdata_axi_m2_o(25)
       , fabric_fpga_rdata_axi_m2_o27                =>  fabric_fpga_rdata_axi_m2_o(26)
       , fabric_fpga_rdata_axi_m2_o28                =>  fabric_fpga_rdata_axi_m2_o(27)
       , fabric_fpga_rdata_axi_m2_o29                =>  fabric_fpga_rdata_axi_m2_o(28)
       , fabric_fpga_rdata_axi_m2_o30                =>  fabric_fpga_rdata_axi_m2_o(29)
       , fabric_fpga_rdata_axi_m2_o31                =>  fabric_fpga_rdata_axi_m2_o(30)
       , fabric_fpga_rdata_axi_m2_o32                =>  fabric_fpga_rdata_axi_m2_o(31)
       , fabric_fpga_rdata_axi_m2_o33                =>  fabric_fpga_rdata_axi_m2_o(32)
       , fabric_fpga_rdata_axi_m2_o34                =>  fabric_fpga_rdata_axi_m2_o(33)
       , fabric_fpga_rdata_axi_m2_o35                =>  fabric_fpga_rdata_axi_m2_o(34)
       , fabric_fpga_rdata_axi_m2_o36                =>  fabric_fpga_rdata_axi_m2_o(35)
       , fabric_fpga_rdata_axi_m2_o37                =>  fabric_fpga_rdata_axi_m2_o(36)
       , fabric_fpga_rdata_axi_m2_o38                =>  fabric_fpga_rdata_axi_m2_o(37)
       , fabric_fpga_rdata_axi_m2_o39                =>  fabric_fpga_rdata_axi_m2_o(38)
       , fabric_fpga_rdata_axi_m2_o40                =>  fabric_fpga_rdata_axi_m2_o(39)
       , fabric_fpga_rdata_axi_m2_o41                =>  fabric_fpga_rdata_axi_m2_o(40)
       , fabric_fpga_rdata_axi_m2_o42                =>  fabric_fpga_rdata_axi_m2_o(41)
       , fabric_fpga_rdata_axi_m2_o43                =>  fabric_fpga_rdata_axi_m2_o(42)
       , fabric_fpga_rdata_axi_m2_o44                =>  fabric_fpga_rdata_axi_m2_o(43)
       , fabric_fpga_rdata_axi_m2_o45                =>  fabric_fpga_rdata_axi_m2_o(44)
       , fabric_fpga_rdata_axi_m2_o46                =>  fabric_fpga_rdata_axi_m2_o(45)
       , fabric_fpga_rdata_axi_m2_o47                =>  fabric_fpga_rdata_axi_m2_o(46)
       , fabric_fpga_rdata_axi_m2_o48                =>  fabric_fpga_rdata_axi_m2_o(47)
       , fabric_fpga_rdata_axi_m2_o49                =>  fabric_fpga_rdata_axi_m2_o(48)
       , fabric_fpga_rdata_axi_m2_o50                =>  fabric_fpga_rdata_axi_m2_o(49)
       , fabric_fpga_rdata_axi_m2_o51                =>  fabric_fpga_rdata_axi_m2_o(50)
       , fabric_fpga_rdata_axi_m2_o52                =>  fabric_fpga_rdata_axi_m2_o(51)
       , fabric_fpga_rdata_axi_m2_o53                =>  fabric_fpga_rdata_axi_m2_o(52)
       , fabric_fpga_rdata_axi_m2_o54                =>  fabric_fpga_rdata_axi_m2_o(53)
       , fabric_fpga_rdata_axi_m2_o55                =>  fabric_fpga_rdata_axi_m2_o(54)
       , fabric_fpga_rdata_axi_m2_o56                =>  fabric_fpga_rdata_axi_m2_o(55)
       , fabric_fpga_rdata_axi_m2_o57                =>  fabric_fpga_rdata_axi_m2_o(56)
       , fabric_fpga_rdata_axi_m2_o58                =>  fabric_fpga_rdata_axi_m2_o(57)
       , fabric_fpga_rdata_axi_m2_o59                =>  fabric_fpga_rdata_axi_m2_o(58)
       , fabric_fpga_rdata_axi_m2_o60                =>  fabric_fpga_rdata_axi_m2_o(59)
       , fabric_fpga_rdata_axi_m2_o61                =>  fabric_fpga_rdata_axi_m2_o(60)
       , fabric_fpga_rdata_axi_m2_o62                =>  fabric_fpga_rdata_axi_m2_o(61)
       , fabric_fpga_rdata_axi_m2_o63                =>  fabric_fpga_rdata_axi_m2_o(62)
       , fabric_fpga_rdata_axi_m2_o64                =>  fabric_fpga_rdata_axi_m2_o(63)
       , fabric_fpga_rdata_axi_m2_o65                =>  fabric_fpga_rdata_axi_m2_o(64)
       , fabric_fpga_rdata_axi_m2_o66                =>  fabric_fpga_rdata_axi_m2_o(65)
       , fabric_fpga_rdata_axi_m2_o67                =>  fabric_fpga_rdata_axi_m2_o(66)
       , fabric_fpga_rdata_axi_m2_o68                =>  fabric_fpga_rdata_axi_m2_o(67)
       , fabric_fpga_rdata_axi_m2_o69                =>  fabric_fpga_rdata_axi_m2_o(68)
       , fabric_fpga_rdata_axi_m2_o70                =>  fabric_fpga_rdata_axi_m2_o(69)
       , fabric_fpga_rdata_axi_m2_o71                =>  fabric_fpga_rdata_axi_m2_o(70)
       , fabric_fpga_rdata_axi_m2_o72                =>  fabric_fpga_rdata_axi_m2_o(71)
       , fabric_fpga_rdata_axi_m2_o73                =>  fabric_fpga_rdata_axi_m2_o(72)
       , fabric_fpga_rdata_axi_m2_o74                =>  fabric_fpga_rdata_axi_m2_o(73)
       , fabric_fpga_rdata_axi_m2_o75                =>  fabric_fpga_rdata_axi_m2_o(74)
       , fabric_fpga_rdata_axi_m2_o76                =>  fabric_fpga_rdata_axi_m2_o(75)
       , fabric_fpga_rdata_axi_m2_o77                =>  fabric_fpga_rdata_axi_m2_o(76)
       , fabric_fpga_rdata_axi_m2_o78                =>  fabric_fpga_rdata_axi_m2_o(77)
       , fabric_fpga_rdata_axi_m2_o79                =>  fabric_fpga_rdata_axi_m2_o(78)
       , fabric_fpga_rdata_axi_m2_o80                =>  fabric_fpga_rdata_axi_m2_o(79)
       , fabric_fpga_rdata_axi_m2_o81                =>  fabric_fpga_rdata_axi_m2_o(80)
       , fabric_fpga_rdata_axi_m2_o82                =>  fabric_fpga_rdata_axi_m2_o(81)
       , fabric_fpga_rdata_axi_m2_o83                =>  fabric_fpga_rdata_axi_m2_o(82)
       , fabric_fpga_rdata_axi_m2_o84                =>  fabric_fpga_rdata_axi_m2_o(83)
       , fabric_fpga_rdata_axi_m2_o85                =>  fabric_fpga_rdata_axi_m2_o(84)
       , fabric_fpga_rdata_axi_m2_o86                =>  fabric_fpga_rdata_axi_m2_o(85)
       , fabric_fpga_rdata_axi_m2_o87                =>  fabric_fpga_rdata_axi_m2_o(86)
       , fabric_fpga_rdata_axi_m2_o88                =>  fabric_fpga_rdata_axi_m2_o(87)
       , fabric_fpga_rdata_axi_m2_o89                =>  fabric_fpga_rdata_axi_m2_o(88)
       , fabric_fpga_rdata_axi_m2_o90                =>  fabric_fpga_rdata_axi_m2_o(89)
       , fabric_fpga_rdata_axi_m2_o91                =>  fabric_fpga_rdata_axi_m2_o(90)
       , fabric_fpga_rdata_axi_m2_o92                =>  fabric_fpga_rdata_axi_m2_o(91)
       , fabric_fpga_rdata_axi_m2_o93                =>  fabric_fpga_rdata_axi_m2_o(92)
       , fabric_fpga_rdata_axi_m2_o94                =>  fabric_fpga_rdata_axi_m2_o(93)
       , fabric_fpga_rdata_axi_m2_o95                =>  fabric_fpga_rdata_axi_m2_o(94)
       , fabric_fpga_rdata_axi_m2_o96                =>  fabric_fpga_rdata_axi_m2_o(95)
       , fabric_fpga_rdata_axi_m2_o97                =>  fabric_fpga_rdata_axi_m2_o(96)
       , fabric_fpga_rdata_axi_m2_o98                =>  fabric_fpga_rdata_axi_m2_o(97)
       , fabric_fpga_rdata_axi_m2_o99                =>  fabric_fpga_rdata_axi_m2_o(98)
       , fabric_fpga_rdata_axi_m2_o100               =>  fabric_fpga_rdata_axi_m2_o(99)
       , fabric_fpga_rdata_axi_m2_o101               =>  fabric_fpga_rdata_axi_m2_o(100)
       , fabric_fpga_rdata_axi_m2_o102               =>  fabric_fpga_rdata_axi_m2_o(101)
       , fabric_fpga_rdata_axi_m2_o103               =>  fabric_fpga_rdata_axi_m2_o(102)
       , fabric_fpga_rdata_axi_m2_o104               =>  fabric_fpga_rdata_axi_m2_o(103)
       , fabric_fpga_rdata_axi_m2_o105               =>  fabric_fpga_rdata_axi_m2_o(104)
       , fabric_fpga_rdata_axi_m2_o106               =>  fabric_fpga_rdata_axi_m2_o(105)
       , fabric_fpga_rdata_axi_m2_o107               =>  fabric_fpga_rdata_axi_m2_o(106)
       , fabric_fpga_rdata_axi_m2_o108               =>  fabric_fpga_rdata_axi_m2_o(107)
       , fabric_fpga_rdata_axi_m2_o109               =>  fabric_fpga_rdata_axi_m2_o(108)
       , fabric_fpga_rdata_axi_m2_o110               =>  fabric_fpga_rdata_axi_m2_o(109)
       , fabric_fpga_rdata_axi_m2_o111               =>  fabric_fpga_rdata_axi_m2_o(110)
       , fabric_fpga_rdata_axi_m2_o112               =>  fabric_fpga_rdata_axi_m2_o(111)
       , fabric_fpga_rdata_axi_m2_o113               =>  fabric_fpga_rdata_axi_m2_o(112)
       , fabric_fpga_rdata_axi_m2_o114               =>  fabric_fpga_rdata_axi_m2_o(113)
       , fabric_fpga_rdata_axi_m2_o115               =>  fabric_fpga_rdata_axi_m2_o(114)
       , fabric_fpga_rdata_axi_m2_o116               =>  fabric_fpga_rdata_axi_m2_o(115)
       , fabric_fpga_rdata_axi_m2_o117               =>  fabric_fpga_rdata_axi_m2_o(116)
       , fabric_fpga_rdata_axi_m2_o118               =>  fabric_fpga_rdata_axi_m2_o(117)
       , fabric_fpga_rdata_axi_m2_o119               =>  fabric_fpga_rdata_axi_m2_o(118)
       , fabric_fpga_rdata_axi_m2_o120               =>  fabric_fpga_rdata_axi_m2_o(119)
       , fabric_fpga_rdata_axi_m2_o121               =>  fabric_fpga_rdata_axi_m2_o(120)
       , fabric_fpga_rdata_axi_m2_o122               =>  fabric_fpga_rdata_axi_m2_o(121)
       , fabric_fpga_rdata_axi_m2_o123               =>  fabric_fpga_rdata_axi_m2_o(122)
       , fabric_fpga_rdata_axi_m2_o124               =>  fabric_fpga_rdata_axi_m2_o(123)
       , fabric_fpga_rdata_axi_m2_o125               =>  fabric_fpga_rdata_axi_m2_o(124)
       , fabric_fpga_rdata_axi_m2_o126               =>  fabric_fpga_rdata_axi_m2_o(125)
       , fabric_fpga_rdata_axi_m2_o127               =>  fabric_fpga_rdata_axi_m2_o(126)
       , fabric_fpga_rdata_axi_m2_o128               =>  fabric_fpga_rdata_axi_m2_o(127)
       , fabric_fpga_rid_axi_m2_o1                   =>  fabric_fpga_rid_axi_m2_o(0)
       , fabric_fpga_rid_axi_m2_o2                   =>  fabric_fpga_rid_axi_m2_o(1)
       , fabric_fpga_rid_axi_m2_o3                   =>  fabric_fpga_rid_axi_m2_o(2)
       , fabric_fpga_rid_axi_m2_o4                   =>  fabric_fpga_rid_axi_m2_o(3)
       , fabric_fpga_rid_axi_m2_o5                   =>  fabric_fpga_rid_axi_m2_o(4)
       , fabric_fpga_rlast_axi_m2_o                  =>  fabric_fpga_rlast_axi_m2_o
       , fabric_fpga_rresp_axi_m2_o1                 =>  fabric_fpga_rresp_axi_m2_o(0)
       , fabric_fpga_rresp_axi_m2_o2                 =>  fabric_fpga_rresp_axi_m2_o(1)
       , fabric_fpga_rvalid_axi_m2_o                 =>  fabric_fpga_rvalid_axi_m2_o
       , fabric_fpga_wready_axi_m2_o                 =>  fabric_fpga_wready_axi_m2_o
       , fabric_fpga_araddr_axi_m2_i1                =>  fabric_fpga_araddr_axi_m2_i(0)
       , fabric_fpga_araddr_axi_m2_i2                =>  fabric_fpga_araddr_axi_m2_i(1)
       , fabric_fpga_araddr_axi_m2_i3                =>  fabric_fpga_araddr_axi_m2_i(2)
       , fabric_fpga_araddr_axi_m2_i4                =>  fabric_fpga_araddr_axi_m2_i(3)
       , fabric_fpga_araddr_axi_m2_i5                =>  fabric_fpga_araddr_axi_m2_i(4)
       , fabric_fpga_araddr_axi_m2_i6                =>  fabric_fpga_araddr_axi_m2_i(5)
       , fabric_fpga_araddr_axi_m2_i7                =>  fabric_fpga_araddr_axi_m2_i(6)
       , fabric_fpga_araddr_axi_m2_i8                =>  fabric_fpga_araddr_axi_m2_i(7)
       , fabric_fpga_araddr_axi_m2_i9                =>  fabric_fpga_araddr_axi_m2_i(8)
       , fabric_fpga_araddr_axi_m2_i10               =>  fabric_fpga_araddr_axi_m2_i(9)
       , fabric_fpga_araddr_axi_m2_i11               =>  fabric_fpga_araddr_axi_m2_i(10)
       , fabric_fpga_araddr_axi_m2_i12               =>  fabric_fpga_araddr_axi_m2_i(11)
       , fabric_fpga_araddr_axi_m2_i13               =>  fabric_fpga_araddr_axi_m2_i(12)
       , fabric_fpga_araddr_axi_m2_i14               =>  fabric_fpga_araddr_axi_m2_i(13)
       , fabric_fpga_araddr_axi_m2_i15               =>  fabric_fpga_araddr_axi_m2_i(14)
       , fabric_fpga_araddr_axi_m2_i16               =>  fabric_fpga_araddr_axi_m2_i(15)
       , fabric_fpga_araddr_axi_m2_i17               =>  fabric_fpga_araddr_axi_m2_i(16)
       , fabric_fpga_araddr_axi_m2_i18               =>  fabric_fpga_araddr_axi_m2_i(17)
       , fabric_fpga_araddr_axi_m2_i19               =>  fabric_fpga_araddr_axi_m2_i(18)
       , fabric_fpga_araddr_axi_m2_i20               =>  fabric_fpga_araddr_axi_m2_i(19)
       , fabric_fpga_araddr_axi_m2_i21               =>  fabric_fpga_araddr_axi_m2_i(20)
       , fabric_fpga_araddr_axi_m2_i22               =>  fabric_fpga_araddr_axi_m2_i(21)
       , fabric_fpga_araddr_axi_m2_i23               =>  fabric_fpga_araddr_axi_m2_i(22)
       , fabric_fpga_araddr_axi_m2_i24               =>  fabric_fpga_araddr_axi_m2_i(23)
       , fabric_fpga_araddr_axi_m2_i25               =>  fabric_fpga_araddr_axi_m2_i(24)
       , fabric_fpga_araddr_axi_m2_i26               =>  fabric_fpga_araddr_axi_m2_i(25)
       , fabric_fpga_araddr_axi_m2_i27               =>  fabric_fpga_araddr_axi_m2_i(26)
       , fabric_fpga_araddr_axi_m2_i28               =>  fabric_fpga_araddr_axi_m2_i(27)
       , fabric_fpga_araddr_axi_m2_i29               =>  fabric_fpga_araddr_axi_m2_i(28)
       , fabric_fpga_araddr_axi_m2_i30               =>  fabric_fpga_araddr_axi_m2_i(29)
       , fabric_fpga_araddr_axi_m2_i31               =>  fabric_fpga_araddr_axi_m2_i(30)
       , fabric_fpga_araddr_axi_m2_i32               =>  fabric_fpga_araddr_axi_m2_i(31)
       , fabric_fpga_araddr_axi_m2_i33               =>  fabric_fpga_araddr_axi_m2_i(32)
       , fabric_fpga_araddr_axi_m2_i34               =>  fabric_fpga_araddr_axi_m2_i(33)
       , fabric_fpga_araddr_axi_m2_i35               =>  fabric_fpga_araddr_axi_m2_i(34)
       , fabric_fpga_araddr_axi_m2_i36               =>  fabric_fpga_araddr_axi_m2_i(35)
       , fabric_fpga_araddr_axi_m2_i37               =>  fabric_fpga_araddr_axi_m2_i(36)
       , fabric_fpga_araddr_axi_m2_i38               =>  fabric_fpga_araddr_axi_m2_i(37)
       , fabric_fpga_araddr_axi_m2_i39               =>  fabric_fpga_araddr_axi_m2_i(38)
       , fabric_fpga_araddr_axi_m2_i40               =>  fabric_fpga_araddr_axi_m2_i(39)
       , fabric_fpga_arburst_axi_m2_i1               =>  fabric_fpga_arburst_axi_m2_i(0)
       , fabric_fpga_arburst_axi_m2_i2               =>  fabric_fpga_arburst_axi_m2_i(1)
       , fabric_fpga_arcache_axi_m2_i1               =>  fabric_fpga_arcache_axi_m2_i(0)
       , fabric_fpga_arcache_axi_m2_i2               =>  fabric_fpga_arcache_axi_m2_i(1)
       , fabric_fpga_arcache_axi_m2_i3               =>  fabric_fpga_arcache_axi_m2_i(2)
       , fabric_fpga_arcache_axi_m2_i4               =>  fabric_fpga_arcache_axi_m2_i(3)
       , fabric_fpga_arid_axi_m2_i1                  =>  fabric_fpga_arid_axi_m2_i(0)
       , fabric_fpga_arid_axi_m2_i2                  =>  fabric_fpga_arid_axi_m2_i(1)
       , fabric_fpga_arid_axi_m2_i3                  =>  fabric_fpga_arid_axi_m2_i(2)
       , fabric_fpga_arid_axi_m2_i4                  =>  fabric_fpga_arid_axi_m2_i(3)
       , fabric_fpga_arid_axi_m2_i5                  =>  fabric_fpga_arid_axi_m2_i(4)
       , fabric_fpga_arlen_axi_m2_i1                 =>  fabric_fpga_arlen_axi_m2_i(0)
       , fabric_fpga_arlen_axi_m2_i2                 =>  fabric_fpga_arlen_axi_m2_i(1)
       , fabric_fpga_arlen_axi_m2_i3                 =>  fabric_fpga_arlen_axi_m2_i(2)
       , fabric_fpga_arlen_axi_m2_i4                 =>  fabric_fpga_arlen_axi_m2_i(3)
       , fabric_fpga_arlen_axi_m2_i5                 =>  fabric_fpga_arlen_axi_m2_i(4)
       , fabric_fpga_arlen_axi_m2_i6                 =>  fabric_fpga_arlen_axi_m2_i(5)
       , fabric_fpga_arlen_axi_m2_i7                 =>  fabric_fpga_arlen_axi_m2_i(6)
       , fabric_fpga_arlen_axi_m2_i8                 =>  fabric_fpga_arlen_axi_m2_i(7)
       , fabric_fpga_arlock_axi_m2_i                 =>  fabric_fpga_arlock_axi_m2_i
       , fabric_fpga_arprot_axi_m2_i1                =>  fabric_fpga_arprot_axi_m2_i(0)
       , fabric_fpga_arprot_axi_m2_i2                =>  fabric_fpga_arprot_axi_m2_i(1)
       , fabric_fpga_arprot_axi_m2_i3                =>  fabric_fpga_arprot_axi_m2_i(2)
       , fabric_fpga_arqos_axi_m2_i1                 =>  fabric_fpga_arqos_axi_m2_i(0)
       , fabric_fpga_arqos_axi_m2_i2                 =>  fabric_fpga_arqos_axi_m2_i(1)
       , fabric_fpga_arqos_axi_m2_i3                 =>  fabric_fpga_arqos_axi_m2_i(2)
       , fabric_fpga_arqos_axi_m2_i4                 =>  fabric_fpga_arqos_axi_m2_i(3)
       , fabric_fpga_arsize_axi_m2_i1                =>  fabric_fpga_arsize_axi_m2_i(0)
       , fabric_fpga_arsize_axi_m2_i2                =>  fabric_fpga_arsize_axi_m2_i(1)
       , fabric_fpga_arsize_axi_m2_i3                =>  fabric_fpga_arsize_axi_m2_i(2)
       , fabric_fpga_arvalid_axi_m2_i                =>  fabric_fpga_arvalid_axi_m2_i
       , fabric_fpga_awaddr_axi_m2_i1                =>  fabric_fpga_awaddr_axi_m2_i(0)
       , fabric_fpga_awaddr_axi_m2_i2                =>  fabric_fpga_awaddr_axi_m2_i(1)
       , fabric_fpga_awaddr_axi_m2_i3                =>  fabric_fpga_awaddr_axi_m2_i(2)
       , fabric_fpga_awaddr_axi_m2_i4                =>  fabric_fpga_awaddr_axi_m2_i(3)
       , fabric_fpga_awaddr_axi_m2_i5                =>  fabric_fpga_awaddr_axi_m2_i(4)
       , fabric_fpga_awaddr_axi_m2_i6                =>  fabric_fpga_awaddr_axi_m2_i(5)
       , fabric_fpga_awaddr_axi_m2_i7                =>  fabric_fpga_awaddr_axi_m2_i(6)
       , fabric_fpga_awaddr_axi_m2_i8                =>  fabric_fpga_awaddr_axi_m2_i(7)
       , fabric_fpga_awaddr_axi_m2_i9                =>  fabric_fpga_awaddr_axi_m2_i(8)
       , fabric_fpga_awaddr_axi_m2_i10               =>  fabric_fpga_awaddr_axi_m2_i(9)
       , fabric_fpga_awaddr_axi_m2_i11               =>  fabric_fpga_awaddr_axi_m2_i(10)
       , fabric_fpga_awaddr_axi_m2_i12               =>  fabric_fpga_awaddr_axi_m2_i(11)
       , fabric_fpga_awaddr_axi_m2_i13               =>  fabric_fpga_awaddr_axi_m2_i(12)
       , fabric_fpga_awaddr_axi_m2_i14               =>  fabric_fpga_awaddr_axi_m2_i(13)
       , fabric_fpga_awaddr_axi_m2_i15               =>  fabric_fpga_awaddr_axi_m2_i(14)
       , fabric_fpga_awaddr_axi_m2_i16               =>  fabric_fpga_awaddr_axi_m2_i(15)
       , fabric_fpga_awaddr_axi_m2_i17               =>  fabric_fpga_awaddr_axi_m2_i(16)
       , fabric_fpga_awaddr_axi_m2_i18               =>  fabric_fpga_awaddr_axi_m2_i(17)
       , fabric_fpga_awaddr_axi_m2_i19               =>  fabric_fpga_awaddr_axi_m2_i(18)
       , fabric_fpga_awaddr_axi_m2_i20               =>  fabric_fpga_awaddr_axi_m2_i(19)
       , fabric_fpga_awaddr_axi_m2_i21               =>  fabric_fpga_awaddr_axi_m2_i(20)
       , fabric_fpga_awaddr_axi_m2_i22               =>  fabric_fpga_awaddr_axi_m2_i(21)
       , fabric_fpga_awaddr_axi_m2_i23               =>  fabric_fpga_awaddr_axi_m2_i(22)
       , fabric_fpga_awaddr_axi_m2_i24               =>  fabric_fpga_awaddr_axi_m2_i(23)
       , fabric_fpga_awaddr_axi_m2_i25               =>  fabric_fpga_awaddr_axi_m2_i(24)
       , fabric_fpga_awaddr_axi_m2_i26               =>  fabric_fpga_awaddr_axi_m2_i(25)
       , fabric_fpga_awaddr_axi_m2_i27               =>  fabric_fpga_awaddr_axi_m2_i(26)
       , fabric_fpga_awaddr_axi_m2_i28               =>  fabric_fpga_awaddr_axi_m2_i(27)
       , fabric_fpga_awaddr_axi_m2_i29               =>  fabric_fpga_awaddr_axi_m2_i(28)
       , fabric_fpga_awaddr_axi_m2_i30               =>  fabric_fpga_awaddr_axi_m2_i(29)
       , fabric_fpga_awaddr_axi_m2_i31               =>  fabric_fpga_awaddr_axi_m2_i(30)
       , fabric_fpga_awaddr_axi_m2_i32               =>  fabric_fpga_awaddr_axi_m2_i(31)
       , fabric_fpga_awaddr_axi_m2_i33               =>  fabric_fpga_awaddr_axi_m2_i(32)
       , fabric_fpga_awaddr_axi_m2_i34               =>  fabric_fpga_awaddr_axi_m2_i(33)
       , fabric_fpga_awaddr_axi_m2_i35               =>  fabric_fpga_awaddr_axi_m2_i(34)
       , fabric_fpga_awaddr_axi_m2_i36               =>  fabric_fpga_awaddr_axi_m2_i(35)
       , fabric_fpga_awaddr_axi_m2_i37               =>  fabric_fpga_awaddr_axi_m2_i(36)
       , fabric_fpga_awaddr_axi_m2_i38               =>  fabric_fpga_awaddr_axi_m2_i(37)
       , fabric_fpga_awaddr_axi_m2_i39               =>  fabric_fpga_awaddr_axi_m2_i(38)
       , fabric_fpga_awaddr_axi_m2_i40               =>  fabric_fpga_awaddr_axi_m2_i(39)
       , fabric_fpga_awburst_axi_m2_i1               =>  fabric_fpga_awburst_axi_m2_i(0)
       , fabric_fpga_awburst_axi_m2_i2               =>  fabric_fpga_awburst_axi_m2_i(1)
       , fabric_fpga_awcache_axi_m2_i1               =>  fabric_fpga_awcache_axi_m2_i(0)
       , fabric_fpga_awcache_axi_m2_i2               =>  fabric_fpga_awcache_axi_m2_i(1)
       , fabric_fpga_awcache_axi_m2_i3               =>  fabric_fpga_awcache_axi_m2_i(2)
       , fabric_fpga_awcache_axi_m2_i4               =>  fabric_fpga_awcache_axi_m2_i(3)
       , fabric_fpga_awid_axi_m2_i1                  =>  fabric_fpga_awid_axi_m2_i(0)
       , fabric_fpga_awid_axi_m2_i2                  =>  fabric_fpga_awid_axi_m2_i(1)
       , fabric_fpga_awid_axi_m2_i3                  =>  fabric_fpga_awid_axi_m2_i(2)
       , fabric_fpga_awid_axi_m2_i4                  =>  fabric_fpga_awid_axi_m2_i(3)
       , fabric_fpga_awid_axi_m2_i5                  =>  fabric_fpga_awid_axi_m2_i(4)
       , fabric_fpga_awlen_axi_m2_i1                 =>  fabric_fpga_awlen_axi_m2_i(0)
       , fabric_fpga_awlen_axi_m2_i2                 =>  fabric_fpga_awlen_axi_m2_i(1)
       , fabric_fpga_awlen_axi_m2_i3                 =>  fabric_fpga_awlen_axi_m2_i(2)
       , fabric_fpga_awlen_axi_m2_i4                 =>  fabric_fpga_awlen_axi_m2_i(3)
       , fabric_fpga_awlen_axi_m2_i5                 =>  fabric_fpga_awlen_axi_m2_i(4)
       , fabric_fpga_awlen_axi_m2_i6                 =>  fabric_fpga_awlen_axi_m2_i(5)
       , fabric_fpga_awlen_axi_m2_i7                 =>  fabric_fpga_awlen_axi_m2_i(6)
       , fabric_fpga_awlen_axi_m2_i8                 =>  fabric_fpga_awlen_axi_m2_i(7)
       , fabric_fpga_awlock_axi_m2_i                 =>  fabric_fpga_awlock_axi_m2_i
       , fabric_fpga_awprot_axi_m2_i1                =>  fabric_fpga_awprot_axi_m2_i(0)
       , fabric_fpga_awprot_axi_m2_i2                =>  fabric_fpga_awprot_axi_m2_i(1)
       , fabric_fpga_awprot_axi_m2_i3                =>  fabric_fpga_awprot_axi_m2_i(2)
       , fabric_fpga_awqos_axi_m2_i1                 =>  fabric_fpga_awqos_axi_m2_i(0)
       , fabric_fpga_awqos_axi_m2_i2                 =>  fabric_fpga_awqos_axi_m2_i(1)
       , fabric_fpga_awqos_axi_m2_i3                 =>  fabric_fpga_awqos_axi_m2_i(2)
       , fabric_fpga_awqos_axi_m2_i4                 =>  fabric_fpga_awqos_axi_m2_i(3)
       , fabric_fpga_awsize_axi_m2_i1                =>  fabric_fpga_awsize_axi_m2_i(0)
       , fabric_fpga_awsize_axi_m2_i2                =>  fabric_fpga_awsize_axi_m2_i(1)
       , fabric_fpga_awsize_axi_m2_i3                =>  fabric_fpga_awsize_axi_m2_i(2)
       , fabric_fpga_awvalid_axi_m2_i                =>  fabric_fpga_awvalid_axi_m2_i
       , fabric_fpga_bready_axi_m2_i                 =>  fabric_fpga_bready_axi_m2_i
       , fabric_fpga_dma_last_m2_i1                  =>  fabric_fpga_dma_last_m2_i(0)
       , fabric_fpga_dma_last_m2_i2                  =>  fabric_fpga_dma_last_m2_i(1)
       , fabric_fpga_dma_last_m2_i3                  =>  fabric_fpga_dma_last_m2_i(2)
       , fabric_fpga_dma_last_m2_i4                  =>  fabric_fpga_dma_last_m2_i(3)
       , fabric_fpga_dma_last_m2_i5                  =>  fabric_fpga_dma_last_m2_i(4)
       , fabric_fpga_dma_last_m2_i6                  =>  fabric_fpga_dma_last_m2_i(5)
       , fabric_fpga_dma_req_m2_i1                   =>  fabric_fpga_dma_req_m2_i(0)
       , fabric_fpga_dma_req_m2_i2                   =>  fabric_fpga_dma_req_m2_i(1)
       , fabric_fpga_dma_req_m2_i3                   =>  fabric_fpga_dma_req_m2_i(2)
       , fabric_fpga_dma_req_m2_i4                   =>  fabric_fpga_dma_req_m2_i(3)
       , fabric_fpga_dma_req_m2_i5                   =>  fabric_fpga_dma_req_m2_i(4)
       , fabric_fpga_dma_req_m2_i6                   =>  fabric_fpga_dma_req_m2_i(5)
       , fabric_fpga_dma_single_m2_i1                =>  fabric_fpga_dma_single_m2_i(0)
       , fabric_fpga_dma_single_m2_i2                =>  fabric_fpga_dma_single_m2_i(1)
       , fabric_fpga_dma_single_m2_i3                =>  fabric_fpga_dma_single_m2_i(2)
       , fabric_fpga_dma_single_m2_i4                =>  fabric_fpga_dma_single_m2_i(3)
       , fabric_fpga_dma_single_m2_i5                =>  fabric_fpga_dma_single_m2_i(4)
       , fabric_fpga_dma_single_m2_i6                =>  fabric_fpga_dma_single_m2_i(5)
       , fabric_fpga_rready_axi_m2_i                 =>  fabric_fpga_rready_axi_m2_i
       , fabric_fpga_wdata_axi_m2_i1                 =>  fabric_fpga_wdata_axi_m2_i(0)
       , fabric_fpga_wdata_axi_m2_i2                 =>  fabric_fpga_wdata_axi_m2_i(1)
       , fabric_fpga_wdata_axi_m2_i3                 =>  fabric_fpga_wdata_axi_m2_i(2)
       , fabric_fpga_wdata_axi_m2_i4                 =>  fabric_fpga_wdata_axi_m2_i(3)
       , fabric_fpga_wdata_axi_m2_i5                 =>  fabric_fpga_wdata_axi_m2_i(4)
       , fabric_fpga_wdata_axi_m2_i6                 =>  fabric_fpga_wdata_axi_m2_i(5)
       , fabric_fpga_wdata_axi_m2_i7                 =>  fabric_fpga_wdata_axi_m2_i(6)
       , fabric_fpga_wdata_axi_m2_i8                 =>  fabric_fpga_wdata_axi_m2_i(7)
       , fabric_fpga_wdata_axi_m2_i9                 =>  fabric_fpga_wdata_axi_m2_i(8)
       , fabric_fpga_wdata_axi_m2_i10                =>  fabric_fpga_wdata_axi_m2_i(9)
       , fabric_fpga_wdata_axi_m2_i11                =>  fabric_fpga_wdata_axi_m2_i(10)
       , fabric_fpga_wdata_axi_m2_i12                =>  fabric_fpga_wdata_axi_m2_i(11)
       , fabric_fpga_wdata_axi_m2_i13                =>  fabric_fpga_wdata_axi_m2_i(12)
       , fabric_fpga_wdata_axi_m2_i14                =>  fabric_fpga_wdata_axi_m2_i(13)
       , fabric_fpga_wdata_axi_m2_i15                =>  fabric_fpga_wdata_axi_m2_i(14)
       , fabric_fpga_wdata_axi_m2_i16                =>  fabric_fpga_wdata_axi_m2_i(15)
       , fabric_fpga_wdata_axi_m2_i17                =>  fabric_fpga_wdata_axi_m2_i(16)
       , fabric_fpga_wdata_axi_m2_i18                =>  fabric_fpga_wdata_axi_m2_i(17)
       , fabric_fpga_wdata_axi_m2_i19                =>  fabric_fpga_wdata_axi_m2_i(18)
       , fabric_fpga_wdata_axi_m2_i20                =>  fabric_fpga_wdata_axi_m2_i(19)
       , fabric_fpga_wdata_axi_m2_i21                =>  fabric_fpga_wdata_axi_m2_i(20)
       , fabric_fpga_wdata_axi_m2_i22                =>  fabric_fpga_wdata_axi_m2_i(21)
       , fabric_fpga_wdata_axi_m2_i23                =>  fabric_fpga_wdata_axi_m2_i(22)
       , fabric_fpga_wdata_axi_m2_i24                =>  fabric_fpga_wdata_axi_m2_i(23)
       , fabric_fpga_wdata_axi_m2_i25                =>  fabric_fpga_wdata_axi_m2_i(24)
       , fabric_fpga_wdata_axi_m2_i26                =>  fabric_fpga_wdata_axi_m2_i(25)
       , fabric_fpga_wdata_axi_m2_i27                =>  fabric_fpga_wdata_axi_m2_i(26)
       , fabric_fpga_wdata_axi_m2_i28                =>  fabric_fpga_wdata_axi_m2_i(27)
       , fabric_fpga_wdata_axi_m2_i29                =>  fabric_fpga_wdata_axi_m2_i(28)
       , fabric_fpga_wdata_axi_m2_i30                =>  fabric_fpga_wdata_axi_m2_i(29)
       , fabric_fpga_wdata_axi_m2_i31                =>  fabric_fpga_wdata_axi_m2_i(30)
       , fabric_fpga_wdata_axi_m2_i32                =>  fabric_fpga_wdata_axi_m2_i(31)
       , fabric_fpga_wdata_axi_m2_i33                =>  fabric_fpga_wdata_axi_m2_i(32)
       , fabric_fpga_wdata_axi_m2_i34                =>  fabric_fpga_wdata_axi_m2_i(33)
       , fabric_fpga_wdata_axi_m2_i35                =>  fabric_fpga_wdata_axi_m2_i(34)
       , fabric_fpga_wdata_axi_m2_i36                =>  fabric_fpga_wdata_axi_m2_i(35)
       , fabric_fpga_wdata_axi_m2_i37                =>  fabric_fpga_wdata_axi_m2_i(36)
       , fabric_fpga_wdata_axi_m2_i38                =>  fabric_fpga_wdata_axi_m2_i(37)
       , fabric_fpga_wdata_axi_m2_i39                =>  fabric_fpga_wdata_axi_m2_i(38)
       , fabric_fpga_wdata_axi_m2_i40                =>  fabric_fpga_wdata_axi_m2_i(39)
       , fabric_fpga_wdata_axi_m2_i41                =>  fabric_fpga_wdata_axi_m2_i(40)
       , fabric_fpga_wdata_axi_m2_i42                =>  fabric_fpga_wdata_axi_m2_i(41)
       , fabric_fpga_wdata_axi_m2_i43                =>  fabric_fpga_wdata_axi_m2_i(42)
       , fabric_fpga_wdata_axi_m2_i44                =>  fabric_fpga_wdata_axi_m2_i(43)
       , fabric_fpga_wdata_axi_m2_i45                =>  fabric_fpga_wdata_axi_m2_i(44)
       , fabric_fpga_wdata_axi_m2_i46                =>  fabric_fpga_wdata_axi_m2_i(45)
       , fabric_fpga_wdata_axi_m2_i47                =>  fabric_fpga_wdata_axi_m2_i(46)
       , fabric_fpga_wdata_axi_m2_i48                =>  fabric_fpga_wdata_axi_m2_i(47)
       , fabric_fpga_wdata_axi_m2_i49                =>  fabric_fpga_wdata_axi_m2_i(48)
       , fabric_fpga_wdata_axi_m2_i50                =>  fabric_fpga_wdata_axi_m2_i(49)
       , fabric_fpga_wdata_axi_m2_i51                =>  fabric_fpga_wdata_axi_m2_i(50)
       , fabric_fpga_wdata_axi_m2_i52                =>  fabric_fpga_wdata_axi_m2_i(51)
       , fabric_fpga_wdata_axi_m2_i53                =>  fabric_fpga_wdata_axi_m2_i(52)
       , fabric_fpga_wdata_axi_m2_i54                =>  fabric_fpga_wdata_axi_m2_i(53)
       , fabric_fpga_wdata_axi_m2_i55                =>  fabric_fpga_wdata_axi_m2_i(54)
       , fabric_fpga_wdata_axi_m2_i56                =>  fabric_fpga_wdata_axi_m2_i(55)
       , fabric_fpga_wdata_axi_m2_i57                =>  fabric_fpga_wdata_axi_m2_i(56)
       , fabric_fpga_wdata_axi_m2_i58                =>  fabric_fpga_wdata_axi_m2_i(57)
       , fabric_fpga_wdata_axi_m2_i59                =>  fabric_fpga_wdata_axi_m2_i(58)
       , fabric_fpga_wdata_axi_m2_i60                =>  fabric_fpga_wdata_axi_m2_i(59)
       , fabric_fpga_wdata_axi_m2_i61                =>  fabric_fpga_wdata_axi_m2_i(60)
       , fabric_fpga_wdata_axi_m2_i62                =>  fabric_fpga_wdata_axi_m2_i(61)
       , fabric_fpga_wdata_axi_m2_i63                =>  fabric_fpga_wdata_axi_m2_i(62)
       , fabric_fpga_wdata_axi_m2_i64                =>  fabric_fpga_wdata_axi_m2_i(63)
       , fabric_fpga_wdata_axi_m2_i65                =>  fabric_fpga_wdata_axi_m2_i(64)
       , fabric_fpga_wdata_axi_m2_i66                =>  fabric_fpga_wdata_axi_m2_i(65)
       , fabric_fpga_wdata_axi_m2_i67                =>  fabric_fpga_wdata_axi_m2_i(66)
       , fabric_fpga_wdata_axi_m2_i68                =>  fabric_fpga_wdata_axi_m2_i(67)
       , fabric_fpga_wdata_axi_m2_i69                =>  fabric_fpga_wdata_axi_m2_i(68)
       , fabric_fpga_wdata_axi_m2_i70                =>  fabric_fpga_wdata_axi_m2_i(69)
       , fabric_fpga_wdata_axi_m2_i71                =>  fabric_fpga_wdata_axi_m2_i(70)
       , fabric_fpga_wdata_axi_m2_i72                =>  fabric_fpga_wdata_axi_m2_i(71)
       , fabric_fpga_wdata_axi_m2_i73                =>  fabric_fpga_wdata_axi_m2_i(72)
       , fabric_fpga_wdata_axi_m2_i74                =>  fabric_fpga_wdata_axi_m2_i(73)
       , fabric_fpga_wdata_axi_m2_i75                =>  fabric_fpga_wdata_axi_m2_i(74)
       , fabric_fpga_wdata_axi_m2_i76                =>  fabric_fpga_wdata_axi_m2_i(75)
       , fabric_fpga_wdata_axi_m2_i77                =>  fabric_fpga_wdata_axi_m2_i(76)
       , fabric_fpga_wdata_axi_m2_i78                =>  fabric_fpga_wdata_axi_m2_i(77)
       , fabric_fpga_wdata_axi_m2_i79                =>  fabric_fpga_wdata_axi_m2_i(78)
       , fabric_fpga_wdata_axi_m2_i80                =>  fabric_fpga_wdata_axi_m2_i(79)
       , fabric_fpga_wdata_axi_m2_i81                =>  fabric_fpga_wdata_axi_m2_i(80)
       , fabric_fpga_wdata_axi_m2_i82                =>  fabric_fpga_wdata_axi_m2_i(81)
       , fabric_fpga_wdata_axi_m2_i83                =>  fabric_fpga_wdata_axi_m2_i(82)
       , fabric_fpga_wdata_axi_m2_i84                =>  fabric_fpga_wdata_axi_m2_i(83)
       , fabric_fpga_wdata_axi_m2_i85                =>  fabric_fpga_wdata_axi_m2_i(84)
       , fabric_fpga_wdata_axi_m2_i86                =>  fabric_fpga_wdata_axi_m2_i(85)
       , fabric_fpga_wdata_axi_m2_i87                =>  fabric_fpga_wdata_axi_m2_i(86)
       , fabric_fpga_wdata_axi_m2_i88                =>  fabric_fpga_wdata_axi_m2_i(87)
       , fabric_fpga_wdata_axi_m2_i89                =>  fabric_fpga_wdata_axi_m2_i(88)
       , fabric_fpga_wdata_axi_m2_i90                =>  fabric_fpga_wdata_axi_m2_i(89)
       , fabric_fpga_wdata_axi_m2_i91                =>  fabric_fpga_wdata_axi_m2_i(90)
       , fabric_fpga_wdata_axi_m2_i92                =>  fabric_fpga_wdata_axi_m2_i(91)
       , fabric_fpga_wdata_axi_m2_i93                =>  fabric_fpga_wdata_axi_m2_i(92)
       , fabric_fpga_wdata_axi_m2_i94                =>  fabric_fpga_wdata_axi_m2_i(93)
       , fabric_fpga_wdata_axi_m2_i95                =>  fabric_fpga_wdata_axi_m2_i(94)
       , fabric_fpga_wdata_axi_m2_i96                =>  fabric_fpga_wdata_axi_m2_i(95)
       , fabric_fpga_wdata_axi_m2_i97                =>  fabric_fpga_wdata_axi_m2_i(96)
       , fabric_fpga_wdata_axi_m2_i98                =>  fabric_fpga_wdata_axi_m2_i(97)
       , fabric_fpga_wdata_axi_m2_i99                =>  fabric_fpga_wdata_axi_m2_i(98)
       , fabric_fpga_wdata_axi_m2_i100               =>  fabric_fpga_wdata_axi_m2_i(99)
       , fabric_fpga_wdata_axi_m2_i101               =>  fabric_fpga_wdata_axi_m2_i(100)
       , fabric_fpga_wdata_axi_m2_i102               =>  fabric_fpga_wdata_axi_m2_i(101)
       , fabric_fpga_wdata_axi_m2_i103               =>  fabric_fpga_wdata_axi_m2_i(102)
       , fabric_fpga_wdata_axi_m2_i104               =>  fabric_fpga_wdata_axi_m2_i(103)
       , fabric_fpga_wdata_axi_m2_i105               =>  fabric_fpga_wdata_axi_m2_i(104)
       , fabric_fpga_wdata_axi_m2_i106               =>  fabric_fpga_wdata_axi_m2_i(105)
       , fabric_fpga_wdata_axi_m2_i107               =>  fabric_fpga_wdata_axi_m2_i(106)
       , fabric_fpga_wdata_axi_m2_i108               =>  fabric_fpga_wdata_axi_m2_i(107)
       , fabric_fpga_wdata_axi_m2_i109               =>  fabric_fpga_wdata_axi_m2_i(108)
       , fabric_fpga_wdata_axi_m2_i110               =>  fabric_fpga_wdata_axi_m2_i(109)
       , fabric_fpga_wdata_axi_m2_i111               =>  fabric_fpga_wdata_axi_m2_i(110)
       , fabric_fpga_wdata_axi_m2_i112               =>  fabric_fpga_wdata_axi_m2_i(111)
       , fabric_fpga_wdata_axi_m2_i113               =>  fabric_fpga_wdata_axi_m2_i(112)
       , fabric_fpga_wdata_axi_m2_i114               =>  fabric_fpga_wdata_axi_m2_i(113)
       , fabric_fpga_wdata_axi_m2_i115               =>  fabric_fpga_wdata_axi_m2_i(114)
       , fabric_fpga_wdata_axi_m2_i116               =>  fabric_fpga_wdata_axi_m2_i(115)
       , fabric_fpga_wdata_axi_m2_i117               =>  fabric_fpga_wdata_axi_m2_i(116)
       , fabric_fpga_wdata_axi_m2_i118               =>  fabric_fpga_wdata_axi_m2_i(117)
       , fabric_fpga_wdata_axi_m2_i119               =>  fabric_fpga_wdata_axi_m2_i(118)
       , fabric_fpga_wdata_axi_m2_i120               =>  fabric_fpga_wdata_axi_m2_i(119)
       , fabric_fpga_wdata_axi_m2_i121               =>  fabric_fpga_wdata_axi_m2_i(120)
       , fabric_fpga_wdata_axi_m2_i122               =>  fabric_fpga_wdata_axi_m2_i(121)
       , fabric_fpga_wdata_axi_m2_i123               =>  fabric_fpga_wdata_axi_m2_i(122)
       , fabric_fpga_wdata_axi_m2_i124               =>  fabric_fpga_wdata_axi_m2_i(123)
       , fabric_fpga_wdata_axi_m2_i125               =>  fabric_fpga_wdata_axi_m2_i(124)
       , fabric_fpga_wdata_axi_m2_i126               =>  fabric_fpga_wdata_axi_m2_i(125)
       , fabric_fpga_wdata_axi_m2_i127               =>  fabric_fpga_wdata_axi_m2_i(126)
       , fabric_fpga_wdata_axi_m2_i128               =>  fabric_fpga_wdata_axi_m2_i(127)
       , fabric_fpga_wlast_axi_m2_i                  =>  fabric_fpga_wlast_axi_m2_i
       , fabric_fpga_wstrb_axi_m2_i1                 =>  fabric_fpga_wstrb_axi_m2_i(0)
       , fabric_fpga_wstrb_axi_m2_i2                 =>  fabric_fpga_wstrb_axi_m2_i(1)
       , fabric_fpga_wstrb_axi_m2_i3                 =>  fabric_fpga_wstrb_axi_m2_i(2)
       , fabric_fpga_wstrb_axi_m2_i4                 =>  fabric_fpga_wstrb_axi_m2_i(3)
       , fabric_fpga_wstrb_axi_m2_i5                 =>  fabric_fpga_wstrb_axi_m2_i(4)
       , fabric_fpga_wstrb_axi_m2_i6                 =>  fabric_fpga_wstrb_axi_m2_i(5)
       , fabric_fpga_wstrb_axi_m2_i7                 =>  fabric_fpga_wstrb_axi_m2_i(6)
       , fabric_fpga_wstrb_axi_m2_i8                 =>  fabric_fpga_wstrb_axi_m2_i(7)
       , fabric_fpga_wstrb_axi_m2_i9                 =>  fabric_fpga_wstrb_axi_m2_i(8)
       , fabric_fpga_wstrb_axi_m2_i10                =>  fabric_fpga_wstrb_axi_m2_i(9)
       , fabric_fpga_wstrb_axi_m2_i11                =>  fabric_fpga_wstrb_axi_m2_i(10)
       , fabric_fpga_wstrb_axi_m2_i12                =>  fabric_fpga_wstrb_axi_m2_i(11)
       , fabric_fpga_wstrb_axi_m2_i13                =>  fabric_fpga_wstrb_axi_m2_i(12)
       , fabric_fpga_wstrb_axi_m2_i14                =>  fabric_fpga_wstrb_axi_m2_i(13)
       , fabric_fpga_wstrb_axi_m2_i15                =>  fabric_fpga_wstrb_axi_m2_i(14)
       , fabric_fpga_wstrb_axi_m2_i16                =>  fabric_fpga_wstrb_axi_m2_i(15)
       , fabric_fpga_wvalid_axi_m2_i                 =>  fabric_fpga_wvalid_axi_m2_i
       , fabric_fpga_ddr0_arready_o                  =>  fabric_fpga_ddr0_arready_o
       , fabric_fpga_ddr0_awready_o                  =>  fabric_fpga_ddr0_awready_o
       , fabric_fpga_ddr0_bid_o1                     =>  fabric_fpga_ddr0_bid_o(0)
       , fabric_fpga_ddr0_bid_o2                     =>  fabric_fpga_ddr0_bid_o(1)
       , fabric_fpga_ddr0_bid_o3                     =>  fabric_fpga_ddr0_bid_o(2)
       , fabric_fpga_ddr0_bid_o4                     =>  fabric_fpga_ddr0_bid_o(3)
       , fabric_fpga_ddr0_bid_o5                     =>  fabric_fpga_ddr0_bid_o(4)
       , fabric_fpga_ddr0_bresp_o1                   =>  fabric_fpga_ddr0_bresp_o(0)
       , fabric_fpga_ddr0_bresp_o2                   =>  fabric_fpga_ddr0_bresp_o(1)
       , fabric_fpga_ddr0_bvalid_o                   =>  fabric_fpga_ddr0_bvalid_o
       , fabric_fpga_ddr0_rdata_o1                   =>  fabric_fpga_ddr0_rdata_o(0)
       , fabric_fpga_ddr0_rdata_o2                   =>  fabric_fpga_ddr0_rdata_o(1)
       , fabric_fpga_ddr0_rdata_o3                   =>  fabric_fpga_ddr0_rdata_o(2)
       , fabric_fpga_ddr0_rdata_o4                   =>  fabric_fpga_ddr0_rdata_o(3)
       , fabric_fpga_ddr0_rdata_o5                   =>  fabric_fpga_ddr0_rdata_o(4)
       , fabric_fpga_ddr0_rdata_o6                   =>  fabric_fpga_ddr0_rdata_o(5)
       , fabric_fpga_ddr0_rdata_o7                   =>  fabric_fpga_ddr0_rdata_o(6)
       , fabric_fpga_ddr0_rdata_o8                   =>  fabric_fpga_ddr0_rdata_o(7)
       , fabric_fpga_ddr0_rdata_o9                   =>  fabric_fpga_ddr0_rdata_o(8)
       , fabric_fpga_ddr0_rdata_o10                  =>  fabric_fpga_ddr0_rdata_o(9)
       , fabric_fpga_ddr0_rdata_o11                  =>  fabric_fpga_ddr0_rdata_o(10)
       , fabric_fpga_ddr0_rdata_o12                  =>  fabric_fpga_ddr0_rdata_o(11)
       , fabric_fpga_ddr0_rdata_o13                  =>  fabric_fpga_ddr0_rdata_o(12)
       , fabric_fpga_ddr0_rdata_o14                  =>  fabric_fpga_ddr0_rdata_o(13)
       , fabric_fpga_ddr0_rdata_o15                  =>  fabric_fpga_ddr0_rdata_o(14)
       , fabric_fpga_ddr0_rdata_o16                  =>  fabric_fpga_ddr0_rdata_o(15)
       , fabric_fpga_ddr0_rdata_o17                  =>  fabric_fpga_ddr0_rdata_o(16)
       , fabric_fpga_ddr0_rdata_o18                  =>  fabric_fpga_ddr0_rdata_o(17)
       , fabric_fpga_ddr0_rdata_o19                  =>  fabric_fpga_ddr0_rdata_o(18)
       , fabric_fpga_ddr0_rdata_o20                  =>  fabric_fpga_ddr0_rdata_o(19)
       , fabric_fpga_ddr0_rdata_o21                  =>  fabric_fpga_ddr0_rdata_o(20)
       , fabric_fpga_ddr0_rdata_o22                  =>  fabric_fpga_ddr0_rdata_o(21)
       , fabric_fpga_ddr0_rdata_o23                  =>  fabric_fpga_ddr0_rdata_o(22)
       , fabric_fpga_ddr0_rdata_o24                  =>  fabric_fpga_ddr0_rdata_o(23)
       , fabric_fpga_ddr0_rdata_o25                  =>  fabric_fpga_ddr0_rdata_o(24)
       , fabric_fpga_ddr0_rdata_o26                  =>  fabric_fpga_ddr0_rdata_o(25)
       , fabric_fpga_ddr0_rdata_o27                  =>  fabric_fpga_ddr0_rdata_o(26)
       , fabric_fpga_ddr0_rdata_o28                  =>  fabric_fpga_ddr0_rdata_o(27)
       , fabric_fpga_ddr0_rdata_o29                  =>  fabric_fpga_ddr0_rdata_o(28)
       , fabric_fpga_ddr0_rdata_o30                  =>  fabric_fpga_ddr0_rdata_o(29)
       , fabric_fpga_ddr0_rdata_o31                  =>  fabric_fpga_ddr0_rdata_o(30)
       , fabric_fpga_ddr0_rdata_o32                  =>  fabric_fpga_ddr0_rdata_o(31)
       , fabric_fpga_ddr0_rdata_o33                  =>  fabric_fpga_ddr0_rdata_o(32)
       , fabric_fpga_ddr0_rdata_o34                  =>  fabric_fpga_ddr0_rdata_o(33)
       , fabric_fpga_ddr0_rdata_o35                  =>  fabric_fpga_ddr0_rdata_o(34)
       , fabric_fpga_ddr0_rdata_o36                  =>  fabric_fpga_ddr0_rdata_o(35)
       , fabric_fpga_ddr0_rdata_o37                  =>  fabric_fpga_ddr0_rdata_o(36)
       , fabric_fpga_ddr0_rdata_o38                  =>  fabric_fpga_ddr0_rdata_o(37)
       , fabric_fpga_ddr0_rdata_o39                  =>  fabric_fpga_ddr0_rdata_o(38)
       , fabric_fpga_ddr0_rdata_o40                  =>  fabric_fpga_ddr0_rdata_o(39)
       , fabric_fpga_ddr0_rdata_o41                  =>  fabric_fpga_ddr0_rdata_o(40)
       , fabric_fpga_ddr0_rdata_o42                  =>  fabric_fpga_ddr0_rdata_o(41)
       , fabric_fpga_ddr0_rdata_o43                  =>  fabric_fpga_ddr0_rdata_o(42)
       , fabric_fpga_ddr0_rdata_o44                  =>  fabric_fpga_ddr0_rdata_o(43)
       , fabric_fpga_ddr0_rdata_o45                  =>  fabric_fpga_ddr0_rdata_o(44)
       , fabric_fpga_ddr0_rdata_o46                  =>  fabric_fpga_ddr0_rdata_o(45)
       , fabric_fpga_ddr0_rdata_o47                  =>  fabric_fpga_ddr0_rdata_o(46)
       , fabric_fpga_ddr0_rdata_o48                  =>  fabric_fpga_ddr0_rdata_o(47)
       , fabric_fpga_ddr0_rdata_o49                  =>  fabric_fpga_ddr0_rdata_o(48)
       , fabric_fpga_ddr0_rdata_o50                  =>  fabric_fpga_ddr0_rdata_o(49)
       , fabric_fpga_ddr0_rdata_o51                  =>  fabric_fpga_ddr0_rdata_o(50)
       , fabric_fpga_ddr0_rdata_o52                  =>  fabric_fpga_ddr0_rdata_o(51)
       , fabric_fpga_ddr0_rdata_o53                  =>  fabric_fpga_ddr0_rdata_o(52)
       , fabric_fpga_ddr0_rdata_o54                  =>  fabric_fpga_ddr0_rdata_o(53)
       , fabric_fpga_ddr0_rdata_o55                  =>  fabric_fpga_ddr0_rdata_o(54)
       , fabric_fpga_ddr0_rdata_o56                  =>  fabric_fpga_ddr0_rdata_o(55)
       , fabric_fpga_ddr0_rdata_o57                  =>  fabric_fpga_ddr0_rdata_o(56)
       , fabric_fpga_ddr0_rdata_o58                  =>  fabric_fpga_ddr0_rdata_o(57)
       , fabric_fpga_ddr0_rdata_o59                  =>  fabric_fpga_ddr0_rdata_o(58)
       , fabric_fpga_ddr0_rdata_o60                  =>  fabric_fpga_ddr0_rdata_o(59)
       , fabric_fpga_ddr0_rdata_o61                  =>  fabric_fpga_ddr0_rdata_o(60)
       , fabric_fpga_ddr0_rdata_o62                  =>  fabric_fpga_ddr0_rdata_o(61)
       , fabric_fpga_ddr0_rdata_o63                  =>  fabric_fpga_ddr0_rdata_o(62)
       , fabric_fpga_ddr0_rdata_o64                  =>  fabric_fpga_ddr0_rdata_o(63)
       , fabric_fpga_ddr0_rdata_o65                  =>  fabric_fpga_ddr0_rdata_o(64)
       , fabric_fpga_ddr0_rdata_o66                  =>  fabric_fpga_ddr0_rdata_o(65)
       , fabric_fpga_ddr0_rdata_o67                  =>  fabric_fpga_ddr0_rdata_o(66)
       , fabric_fpga_ddr0_rdata_o68                  =>  fabric_fpga_ddr0_rdata_o(67)
       , fabric_fpga_ddr0_rdata_o69                  =>  fabric_fpga_ddr0_rdata_o(68)
       , fabric_fpga_ddr0_rdata_o70                  =>  fabric_fpga_ddr0_rdata_o(69)
       , fabric_fpga_ddr0_rdata_o71                  =>  fabric_fpga_ddr0_rdata_o(70)
       , fabric_fpga_ddr0_rdata_o72                  =>  fabric_fpga_ddr0_rdata_o(71)
       , fabric_fpga_ddr0_rdata_o73                  =>  fabric_fpga_ddr0_rdata_o(72)
       , fabric_fpga_ddr0_rdata_o74                  =>  fabric_fpga_ddr0_rdata_o(73)
       , fabric_fpga_ddr0_rdata_o75                  =>  fabric_fpga_ddr0_rdata_o(74)
       , fabric_fpga_ddr0_rdata_o76                  =>  fabric_fpga_ddr0_rdata_o(75)
       , fabric_fpga_ddr0_rdata_o77                  =>  fabric_fpga_ddr0_rdata_o(76)
       , fabric_fpga_ddr0_rdata_o78                  =>  fabric_fpga_ddr0_rdata_o(77)
       , fabric_fpga_ddr0_rdata_o79                  =>  fabric_fpga_ddr0_rdata_o(78)
       , fabric_fpga_ddr0_rdata_o80                  =>  fabric_fpga_ddr0_rdata_o(79)
       , fabric_fpga_ddr0_rdata_o81                  =>  fabric_fpga_ddr0_rdata_o(80)
       , fabric_fpga_ddr0_rdata_o82                  =>  fabric_fpga_ddr0_rdata_o(81)
       , fabric_fpga_ddr0_rdata_o83                  =>  fabric_fpga_ddr0_rdata_o(82)
       , fabric_fpga_ddr0_rdata_o84                  =>  fabric_fpga_ddr0_rdata_o(83)
       , fabric_fpga_ddr0_rdata_o85                  =>  fabric_fpga_ddr0_rdata_o(84)
       , fabric_fpga_ddr0_rdata_o86                  =>  fabric_fpga_ddr0_rdata_o(85)
       , fabric_fpga_ddr0_rdata_o87                  =>  fabric_fpga_ddr0_rdata_o(86)
       , fabric_fpga_ddr0_rdata_o88                  =>  fabric_fpga_ddr0_rdata_o(87)
       , fabric_fpga_ddr0_rdata_o89                  =>  fabric_fpga_ddr0_rdata_o(88)
       , fabric_fpga_ddr0_rdata_o90                  =>  fabric_fpga_ddr0_rdata_o(89)
       , fabric_fpga_ddr0_rdata_o91                  =>  fabric_fpga_ddr0_rdata_o(90)
       , fabric_fpga_ddr0_rdata_o92                  =>  fabric_fpga_ddr0_rdata_o(91)
       , fabric_fpga_ddr0_rdata_o93                  =>  fabric_fpga_ddr0_rdata_o(92)
       , fabric_fpga_ddr0_rdata_o94                  =>  fabric_fpga_ddr0_rdata_o(93)
       , fabric_fpga_ddr0_rdata_o95                  =>  fabric_fpga_ddr0_rdata_o(94)
       , fabric_fpga_ddr0_rdata_o96                  =>  fabric_fpga_ddr0_rdata_o(95)
       , fabric_fpga_ddr0_rdata_o97                  =>  fabric_fpga_ddr0_rdata_o(96)
       , fabric_fpga_ddr0_rdata_o98                  =>  fabric_fpga_ddr0_rdata_o(97)
       , fabric_fpga_ddr0_rdata_o99                  =>  fabric_fpga_ddr0_rdata_o(98)
       , fabric_fpga_ddr0_rdata_o100                 =>  fabric_fpga_ddr0_rdata_o(99)
       , fabric_fpga_ddr0_rdata_o101                 =>  fabric_fpga_ddr0_rdata_o(100)
       , fabric_fpga_ddr0_rdata_o102                 =>  fabric_fpga_ddr0_rdata_o(101)
       , fabric_fpga_ddr0_rdata_o103                 =>  fabric_fpga_ddr0_rdata_o(102)
       , fabric_fpga_ddr0_rdata_o104                 =>  fabric_fpga_ddr0_rdata_o(103)
       , fabric_fpga_ddr0_rdata_o105                 =>  fabric_fpga_ddr0_rdata_o(104)
       , fabric_fpga_ddr0_rdata_o106                 =>  fabric_fpga_ddr0_rdata_o(105)
       , fabric_fpga_ddr0_rdata_o107                 =>  fabric_fpga_ddr0_rdata_o(106)
       , fabric_fpga_ddr0_rdata_o108                 =>  fabric_fpga_ddr0_rdata_o(107)
       , fabric_fpga_ddr0_rdata_o109                 =>  fabric_fpga_ddr0_rdata_o(108)
       , fabric_fpga_ddr0_rdata_o110                 =>  fabric_fpga_ddr0_rdata_o(109)
       , fabric_fpga_ddr0_rdata_o111                 =>  fabric_fpga_ddr0_rdata_o(110)
       , fabric_fpga_ddr0_rdata_o112                 =>  fabric_fpga_ddr0_rdata_o(111)
       , fabric_fpga_ddr0_rdata_o113                 =>  fabric_fpga_ddr0_rdata_o(112)
       , fabric_fpga_ddr0_rdata_o114                 =>  fabric_fpga_ddr0_rdata_o(113)
       , fabric_fpga_ddr0_rdata_o115                 =>  fabric_fpga_ddr0_rdata_o(114)
       , fabric_fpga_ddr0_rdata_o116                 =>  fabric_fpga_ddr0_rdata_o(115)
       , fabric_fpga_ddr0_rdata_o117                 =>  fabric_fpga_ddr0_rdata_o(116)
       , fabric_fpga_ddr0_rdata_o118                 =>  fabric_fpga_ddr0_rdata_o(117)
       , fabric_fpga_ddr0_rdata_o119                 =>  fabric_fpga_ddr0_rdata_o(118)
       , fabric_fpga_ddr0_rdata_o120                 =>  fabric_fpga_ddr0_rdata_o(119)
       , fabric_fpga_ddr0_rdata_o121                 =>  fabric_fpga_ddr0_rdata_o(120)
       , fabric_fpga_ddr0_rdata_o122                 =>  fabric_fpga_ddr0_rdata_o(121)
       , fabric_fpga_ddr0_rdata_o123                 =>  fabric_fpga_ddr0_rdata_o(122)
       , fabric_fpga_ddr0_rdata_o124                 =>  fabric_fpga_ddr0_rdata_o(123)
       , fabric_fpga_ddr0_rdata_o125                 =>  fabric_fpga_ddr0_rdata_o(124)
       , fabric_fpga_ddr0_rdata_o126                 =>  fabric_fpga_ddr0_rdata_o(125)
       , fabric_fpga_ddr0_rdata_o127                 =>  fabric_fpga_ddr0_rdata_o(126)
       , fabric_fpga_ddr0_rdata_o128                 =>  fabric_fpga_ddr0_rdata_o(127)
       , fabric_fpga_ddr0_rid_o1                     =>  fabric_fpga_ddr0_rid_o(0)
       , fabric_fpga_ddr0_rid_o2                     =>  fabric_fpga_ddr0_rid_o(1)
       , fabric_fpga_ddr0_rid_o3                     =>  fabric_fpga_ddr0_rid_o(2)
       , fabric_fpga_ddr0_rid_o4                     =>  fabric_fpga_ddr0_rid_o(3)
       , fabric_fpga_ddr0_rid_o5                     =>  fabric_fpga_ddr0_rid_o(4)
       , fabric_fpga_ddr0_rlast_o                    =>  fabric_fpga_ddr0_rlast_o
       , fabric_fpga_ddr0_rresp_o1                   =>  fabric_fpga_ddr0_rresp_o(0)
       , fabric_fpga_ddr0_rresp_o2                   =>  fabric_fpga_ddr0_rresp_o(1)
       , fabric_fpga_ddr0_rvalid_o                   =>  fabric_fpga_ddr0_rvalid_o
       , fabric_fpga_ddr0_wready_o                   =>  fabric_fpga_ddr0_wready_o
       , fabric_fpga_ddr0_araddr_i1                  =>  fabric_fpga_ddr0_araddr_i(0)
       , fabric_fpga_ddr0_araddr_i2                  =>  fabric_fpga_ddr0_araddr_i(1)
       , fabric_fpga_ddr0_araddr_i3                  =>  fabric_fpga_ddr0_araddr_i(2)
       , fabric_fpga_ddr0_araddr_i4                  =>  fabric_fpga_ddr0_araddr_i(3)
       , fabric_fpga_ddr0_araddr_i5                  =>  fabric_fpga_ddr0_araddr_i(4)
       , fabric_fpga_ddr0_araddr_i6                  =>  fabric_fpga_ddr0_araddr_i(5)
       , fabric_fpga_ddr0_araddr_i7                  =>  fabric_fpga_ddr0_araddr_i(6)
       , fabric_fpga_ddr0_araddr_i8                  =>  fabric_fpga_ddr0_araddr_i(7)
       , fabric_fpga_ddr0_araddr_i9                  =>  fabric_fpga_ddr0_araddr_i(8)
       , fabric_fpga_ddr0_araddr_i10                 =>  fabric_fpga_ddr0_araddr_i(9)
       , fabric_fpga_ddr0_araddr_i11                 =>  fabric_fpga_ddr0_araddr_i(10)
       , fabric_fpga_ddr0_araddr_i12                 =>  fabric_fpga_ddr0_araddr_i(11)
       , fabric_fpga_ddr0_araddr_i13                 =>  fabric_fpga_ddr0_araddr_i(12)
       , fabric_fpga_ddr0_araddr_i14                 =>  fabric_fpga_ddr0_araddr_i(13)
       , fabric_fpga_ddr0_araddr_i15                 =>  fabric_fpga_ddr0_araddr_i(14)
       , fabric_fpga_ddr0_araddr_i16                 =>  fabric_fpga_ddr0_araddr_i(15)
       , fabric_fpga_ddr0_araddr_i17                 =>  fabric_fpga_ddr0_araddr_i(16)
       , fabric_fpga_ddr0_araddr_i18                 =>  fabric_fpga_ddr0_araddr_i(17)
       , fabric_fpga_ddr0_araddr_i19                 =>  fabric_fpga_ddr0_araddr_i(18)
       , fabric_fpga_ddr0_araddr_i20                 =>  fabric_fpga_ddr0_araddr_i(19)
       , fabric_fpga_ddr0_araddr_i21                 =>  fabric_fpga_ddr0_araddr_i(20)
       , fabric_fpga_ddr0_araddr_i22                 =>  fabric_fpga_ddr0_araddr_i(21)
       , fabric_fpga_ddr0_araddr_i23                 =>  fabric_fpga_ddr0_araddr_i(22)
       , fabric_fpga_ddr0_araddr_i24                 =>  fabric_fpga_ddr0_araddr_i(23)
       , fabric_fpga_ddr0_araddr_i25                 =>  fabric_fpga_ddr0_araddr_i(24)
       , fabric_fpga_ddr0_araddr_i26                 =>  fabric_fpga_ddr0_araddr_i(25)
       , fabric_fpga_ddr0_araddr_i27                 =>  fabric_fpga_ddr0_araddr_i(26)
       , fabric_fpga_ddr0_araddr_i28                 =>  fabric_fpga_ddr0_araddr_i(27)
       , fabric_fpga_ddr0_araddr_i29                 =>  fabric_fpga_ddr0_araddr_i(28)
       , fabric_fpga_ddr0_araddr_i30                 =>  fabric_fpga_ddr0_araddr_i(29)
       , fabric_fpga_ddr0_araddr_i31                 =>  fabric_fpga_ddr0_araddr_i(30)
       , fabric_fpga_ddr0_araddr_i32                 =>  fabric_fpga_ddr0_araddr_i(31)
       , fabric_fpga_ddr0_araddr_i33                 =>  fabric_fpga_ddr0_araddr_i(32)
       , fabric_fpga_ddr0_araddr_i34                 =>  fabric_fpga_ddr0_araddr_i(33)
       , fabric_fpga_ddr0_araddr_i35                 =>  fabric_fpga_ddr0_araddr_i(34)
       , fabric_fpga_ddr0_araddr_i36                 =>  fabric_fpga_ddr0_araddr_i(35)
       , fabric_fpga_ddr0_araddr_i37                 =>  fabric_fpga_ddr0_araddr_i(36)
       , fabric_fpga_ddr0_araddr_i38                 =>  fabric_fpga_ddr0_araddr_i(37)
       , fabric_fpga_ddr0_araddr_i39                 =>  fabric_fpga_ddr0_araddr_i(38)
       , fabric_fpga_ddr0_araddr_i40                 =>  fabric_fpga_ddr0_araddr_i(39)
       , fabric_fpga_ddr0_arburst_i1                 =>  fabric_fpga_ddr0_arburst_i(0)
       , fabric_fpga_ddr0_arburst_i2                 =>  fabric_fpga_ddr0_arburst_i(1)
       , fabric_fpga_ddr0_arcache_i1                 =>  fabric_fpga_ddr0_arcache_i(0)
       , fabric_fpga_ddr0_arcache_i2                 =>  fabric_fpga_ddr0_arcache_i(1)
       , fabric_fpga_ddr0_arcache_i3                 =>  fabric_fpga_ddr0_arcache_i(2)
       , fabric_fpga_ddr0_arcache_i4                 =>  fabric_fpga_ddr0_arcache_i(3)
       , fabric_fpga_ddr0_arid_i1                    =>  fabric_fpga_ddr0_arid_i(0)
       , fabric_fpga_ddr0_arid_i2                    =>  fabric_fpga_ddr0_arid_i(1)
       , fabric_fpga_ddr0_arid_i3                    =>  fabric_fpga_ddr0_arid_i(2)
       , fabric_fpga_ddr0_arid_i4                    =>  fabric_fpga_ddr0_arid_i(3)
       , fabric_fpga_ddr0_arid_i5                    =>  fabric_fpga_ddr0_arid_i(4)
       , fabric_fpga_ddr0_arlen_i1                   =>  fabric_fpga_ddr0_arlen_i(0)
       , fabric_fpga_ddr0_arlen_i2                   =>  fabric_fpga_ddr0_arlen_i(1)
       , fabric_fpga_ddr0_arlen_i3                   =>  fabric_fpga_ddr0_arlen_i(2)
       , fabric_fpga_ddr0_arlen_i4                   =>  fabric_fpga_ddr0_arlen_i(3)
       , fabric_fpga_ddr0_arlen_i5                   =>  fabric_fpga_ddr0_arlen_i(4)
       , fabric_fpga_ddr0_arlen_i6                   =>  fabric_fpga_ddr0_arlen_i(5)
       , fabric_fpga_ddr0_arlen_i7                   =>  fabric_fpga_ddr0_arlen_i(6)
       , fabric_fpga_ddr0_arlen_i8                   =>  fabric_fpga_ddr0_arlen_i(7)
       , fabric_fpga_ddr0_arlock_i                   =>  fabric_fpga_ddr0_arlock_i
       , fabric_fpga_ddr0_arprot_i1                  =>  fabric_fpga_ddr0_arprot_i(0)
       , fabric_fpga_ddr0_arprot_i2                  =>  fabric_fpga_ddr0_arprot_i(1)
       , fabric_fpga_ddr0_arprot_i3                  =>  fabric_fpga_ddr0_arprot_i(2)
       , fabric_fpga_ddr0_arqos_i1                   =>  fabric_fpga_ddr0_arqos_i(0)
       , fabric_fpga_ddr0_arqos_i2                   =>  fabric_fpga_ddr0_arqos_i(1)
       , fabric_fpga_ddr0_arqos_i3                   =>  fabric_fpga_ddr0_arqos_i(2)
       , fabric_fpga_ddr0_arqos_i4                   =>  fabric_fpga_ddr0_arqos_i(3)
       , fabric_fpga_ddr0_arsize_i1                  =>  fabric_fpga_ddr0_arsize_i(0)
       , fabric_fpga_ddr0_arsize_i2                  =>  fabric_fpga_ddr0_arsize_i(1)
       , fabric_fpga_ddr0_arsize_i3                  =>  fabric_fpga_ddr0_arsize_i(2)
       , fabric_fpga_ddr0_arvalid_i                  =>  fabric_fpga_ddr0_arvalid_i
       , fabric_fpga_ddr0_awaddr_i1                  =>  fabric_fpga_ddr0_awaddr_i(0)
       , fabric_fpga_ddr0_awaddr_i2                  =>  fabric_fpga_ddr0_awaddr_i(1)
       , fabric_fpga_ddr0_awaddr_i3                  =>  fabric_fpga_ddr0_awaddr_i(2)
       , fabric_fpga_ddr0_awaddr_i4                  =>  fabric_fpga_ddr0_awaddr_i(3)
       , fabric_fpga_ddr0_awaddr_i5                  =>  fabric_fpga_ddr0_awaddr_i(4)
       , fabric_fpga_ddr0_awaddr_i6                  =>  fabric_fpga_ddr0_awaddr_i(5)
       , fabric_fpga_ddr0_awaddr_i7                  =>  fabric_fpga_ddr0_awaddr_i(6)
       , fabric_fpga_ddr0_awaddr_i8                  =>  fabric_fpga_ddr0_awaddr_i(7)
       , fabric_fpga_ddr0_awaddr_i9                  =>  fabric_fpga_ddr0_awaddr_i(8)
       , fabric_fpga_ddr0_awaddr_i10                 =>  fabric_fpga_ddr0_awaddr_i(9)
       , fabric_fpga_ddr0_awaddr_i11                 =>  fabric_fpga_ddr0_awaddr_i(10)
       , fabric_fpga_ddr0_awaddr_i12                 =>  fabric_fpga_ddr0_awaddr_i(11)
       , fabric_fpga_ddr0_awaddr_i13                 =>  fabric_fpga_ddr0_awaddr_i(12)
       , fabric_fpga_ddr0_awaddr_i14                 =>  fabric_fpga_ddr0_awaddr_i(13)
       , fabric_fpga_ddr0_awaddr_i15                 =>  fabric_fpga_ddr0_awaddr_i(14)
       , fabric_fpga_ddr0_awaddr_i16                 =>  fabric_fpga_ddr0_awaddr_i(15)
       , fabric_fpga_ddr0_awaddr_i17                 =>  fabric_fpga_ddr0_awaddr_i(16)
       , fabric_fpga_ddr0_awaddr_i18                 =>  fabric_fpga_ddr0_awaddr_i(17)
       , fabric_fpga_ddr0_awaddr_i19                 =>  fabric_fpga_ddr0_awaddr_i(18)
       , fabric_fpga_ddr0_awaddr_i20                 =>  fabric_fpga_ddr0_awaddr_i(19)
       , fabric_fpga_ddr0_awaddr_i21                 =>  fabric_fpga_ddr0_awaddr_i(20)
       , fabric_fpga_ddr0_awaddr_i22                 =>  fabric_fpga_ddr0_awaddr_i(21)
       , fabric_fpga_ddr0_awaddr_i23                 =>  fabric_fpga_ddr0_awaddr_i(22)
       , fabric_fpga_ddr0_awaddr_i24                 =>  fabric_fpga_ddr0_awaddr_i(23)
       , fabric_fpga_ddr0_awaddr_i25                 =>  fabric_fpga_ddr0_awaddr_i(24)
       , fabric_fpga_ddr0_awaddr_i26                 =>  fabric_fpga_ddr0_awaddr_i(25)
       , fabric_fpga_ddr0_awaddr_i27                 =>  fabric_fpga_ddr0_awaddr_i(26)
       , fabric_fpga_ddr0_awaddr_i28                 =>  fabric_fpga_ddr0_awaddr_i(27)
       , fabric_fpga_ddr0_awaddr_i29                 =>  fabric_fpga_ddr0_awaddr_i(28)
       , fabric_fpga_ddr0_awaddr_i30                 =>  fabric_fpga_ddr0_awaddr_i(29)
       , fabric_fpga_ddr0_awaddr_i31                 =>  fabric_fpga_ddr0_awaddr_i(30)
       , fabric_fpga_ddr0_awaddr_i32                 =>  fabric_fpga_ddr0_awaddr_i(31)
       , fabric_fpga_ddr0_awaddr_i33                 =>  fabric_fpga_ddr0_awaddr_i(32)
       , fabric_fpga_ddr0_awaddr_i34                 =>  fabric_fpga_ddr0_awaddr_i(33)
       , fabric_fpga_ddr0_awaddr_i35                 =>  fabric_fpga_ddr0_awaddr_i(34)
       , fabric_fpga_ddr0_awaddr_i36                 =>  fabric_fpga_ddr0_awaddr_i(35)
       , fabric_fpga_ddr0_awaddr_i37                 =>  fabric_fpga_ddr0_awaddr_i(36)
       , fabric_fpga_ddr0_awaddr_i38                 =>  fabric_fpga_ddr0_awaddr_i(37)
       , fabric_fpga_ddr0_awaddr_i39                 =>  fabric_fpga_ddr0_awaddr_i(38)
       , fabric_fpga_ddr0_awaddr_i40                 =>  fabric_fpga_ddr0_awaddr_i(39)
       , fabric_fpga_ddr0_awburst_i1                 =>  fabric_fpga_ddr0_awburst_i(0)
       , fabric_fpga_ddr0_awburst_i2                 =>  fabric_fpga_ddr0_awburst_i(1)
       , fabric_fpga_ddr0_awcache_i1                 =>  fabric_fpga_ddr0_awcache_i(0)
       , fabric_fpga_ddr0_awcache_i2                 =>  fabric_fpga_ddr0_awcache_i(1)
       , fabric_fpga_ddr0_awcache_i3                 =>  fabric_fpga_ddr0_awcache_i(2)
       , fabric_fpga_ddr0_awcache_i4                 =>  fabric_fpga_ddr0_awcache_i(3)
       , fabric_fpga_ddr0_awid_i1                    =>  fabric_fpga_ddr0_awid_i(0)
       , fabric_fpga_ddr0_awid_i2                    =>  fabric_fpga_ddr0_awid_i(1)
       , fabric_fpga_ddr0_awid_i3                    =>  fabric_fpga_ddr0_awid_i(2)
       , fabric_fpga_ddr0_awid_i4                    =>  fabric_fpga_ddr0_awid_i(3)
       , fabric_fpga_ddr0_awid_i5                    =>  fabric_fpga_ddr0_awid_i(4)
       , fabric_fpga_ddr0_awlen_i1                   =>  fabric_fpga_ddr0_awlen_i(0)
       , fabric_fpga_ddr0_awlen_i2                   =>  fabric_fpga_ddr0_awlen_i(1)
       , fabric_fpga_ddr0_awlen_i3                   =>  fabric_fpga_ddr0_awlen_i(2)
       , fabric_fpga_ddr0_awlen_i4                   =>  fabric_fpga_ddr0_awlen_i(3)
       , fabric_fpga_ddr0_awlen_i5                   =>  fabric_fpga_ddr0_awlen_i(4)
       , fabric_fpga_ddr0_awlen_i6                   =>  fabric_fpga_ddr0_awlen_i(5)
       , fabric_fpga_ddr0_awlen_i7                   =>  fabric_fpga_ddr0_awlen_i(6)
       , fabric_fpga_ddr0_awlen_i8                   =>  fabric_fpga_ddr0_awlen_i(7)
       , fabric_fpga_ddr0_awlock_i                   =>  fabric_fpga_ddr0_awlock_i
       , fabric_fpga_ddr0_awprot_i1                  =>  fabric_fpga_ddr0_awprot_i(0)
       , fabric_fpga_ddr0_awprot_i2                  =>  fabric_fpga_ddr0_awprot_i(1)
       , fabric_fpga_ddr0_awprot_i3                  =>  fabric_fpga_ddr0_awprot_i(2)
       , fabric_fpga_ddr0_awqos_i1                   =>  fabric_fpga_ddr0_awqos_i(0)
       , fabric_fpga_ddr0_awqos_i2                   =>  fabric_fpga_ddr0_awqos_i(1)
       , fabric_fpga_ddr0_awqos_i3                   =>  fabric_fpga_ddr0_awqos_i(2)
       , fabric_fpga_ddr0_awqos_i4                   =>  fabric_fpga_ddr0_awqos_i(3)
       , fabric_fpga_ddr0_awsize_i1                  =>  fabric_fpga_ddr0_awsize_i(0)
       , fabric_fpga_ddr0_awsize_i2                  =>  fabric_fpga_ddr0_awsize_i(1)
       , fabric_fpga_ddr0_awsize_i3                  =>  fabric_fpga_ddr0_awsize_i(2)
       , fabric_fpga_ddr0_awvalid_i                  =>  fabric_fpga_ddr0_awvalid_i
       , fabric_fpga_ddr0_bready_i                   =>  fabric_fpga_ddr0_bready_i
       , fabric_fpga_ddr0_rready_i                   =>  fabric_fpga_ddr0_rready_i
       , fabric_fpga_ddr0_wdata_i1                   =>  fabric_fpga_ddr0_wdata_i(0)
       , fabric_fpga_ddr0_wdata_i2                   =>  fabric_fpga_ddr0_wdata_i(1)
       , fabric_fpga_ddr0_wdata_i3                   =>  fabric_fpga_ddr0_wdata_i(2)
       , fabric_fpga_ddr0_wdata_i4                   =>  fabric_fpga_ddr0_wdata_i(3)
       , fabric_fpga_ddr0_wdata_i5                   =>  fabric_fpga_ddr0_wdata_i(4)
       , fabric_fpga_ddr0_wdata_i6                   =>  fabric_fpga_ddr0_wdata_i(5)
       , fabric_fpga_ddr0_wdata_i7                   =>  fabric_fpga_ddr0_wdata_i(6)
       , fabric_fpga_ddr0_wdata_i8                   =>  fabric_fpga_ddr0_wdata_i(7)
       , fabric_fpga_ddr0_wdata_i9                   =>  fabric_fpga_ddr0_wdata_i(8)
       , fabric_fpga_ddr0_wdata_i10                  =>  fabric_fpga_ddr0_wdata_i(9)
       , fabric_fpga_ddr0_wdata_i11                  =>  fabric_fpga_ddr0_wdata_i(10)
       , fabric_fpga_ddr0_wdata_i12                  =>  fabric_fpga_ddr0_wdata_i(11)
       , fabric_fpga_ddr0_wdata_i13                  =>  fabric_fpga_ddr0_wdata_i(12)
       , fabric_fpga_ddr0_wdata_i14                  =>  fabric_fpga_ddr0_wdata_i(13)
       , fabric_fpga_ddr0_wdata_i15                  =>  fabric_fpga_ddr0_wdata_i(14)
       , fabric_fpga_ddr0_wdata_i16                  =>  fabric_fpga_ddr0_wdata_i(15)
       , fabric_fpga_ddr0_wdata_i17                  =>  fabric_fpga_ddr0_wdata_i(16)
       , fabric_fpga_ddr0_wdata_i18                  =>  fabric_fpga_ddr0_wdata_i(17)
       , fabric_fpga_ddr0_wdata_i19                  =>  fabric_fpga_ddr0_wdata_i(18)
       , fabric_fpga_ddr0_wdata_i20                  =>  fabric_fpga_ddr0_wdata_i(19)
       , fabric_fpga_ddr0_wdata_i21                  =>  fabric_fpga_ddr0_wdata_i(20)
       , fabric_fpga_ddr0_wdata_i22                  =>  fabric_fpga_ddr0_wdata_i(21)
       , fabric_fpga_ddr0_wdata_i23                  =>  fabric_fpga_ddr0_wdata_i(22)
       , fabric_fpga_ddr0_wdata_i24                  =>  fabric_fpga_ddr0_wdata_i(23)
       , fabric_fpga_ddr0_wdata_i25                  =>  fabric_fpga_ddr0_wdata_i(24)
       , fabric_fpga_ddr0_wdata_i26                  =>  fabric_fpga_ddr0_wdata_i(25)
       , fabric_fpga_ddr0_wdata_i27                  =>  fabric_fpga_ddr0_wdata_i(26)
       , fabric_fpga_ddr0_wdata_i28                  =>  fabric_fpga_ddr0_wdata_i(27)
       , fabric_fpga_ddr0_wdata_i29                  =>  fabric_fpga_ddr0_wdata_i(28)
       , fabric_fpga_ddr0_wdata_i30                  =>  fabric_fpga_ddr0_wdata_i(29)
       , fabric_fpga_ddr0_wdata_i31                  =>  fabric_fpga_ddr0_wdata_i(30)
       , fabric_fpga_ddr0_wdata_i32                  =>  fabric_fpga_ddr0_wdata_i(31)
       , fabric_fpga_ddr0_wdata_i33                  =>  fabric_fpga_ddr0_wdata_i(32)
       , fabric_fpga_ddr0_wdata_i34                  =>  fabric_fpga_ddr0_wdata_i(33)
       , fabric_fpga_ddr0_wdata_i35                  =>  fabric_fpga_ddr0_wdata_i(34)
       , fabric_fpga_ddr0_wdata_i36                  =>  fabric_fpga_ddr0_wdata_i(35)
       , fabric_fpga_ddr0_wdata_i37                  =>  fabric_fpga_ddr0_wdata_i(36)
       , fabric_fpga_ddr0_wdata_i38                  =>  fabric_fpga_ddr0_wdata_i(37)
       , fabric_fpga_ddr0_wdata_i39                  =>  fabric_fpga_ddr0_wdata_i(38)
       , fabric_fpga_ddr0_wdata_i40                  =>  fabric_fpga_ddr0_wdata_i(39)
       , fabric_fpga_ddr0_wdata_i41                  =>  fabric_fpga_ddr0_wdata_i(40)
       , fabric_fpga_ddr0_wdata_i42                  =>  fabric_fpga_ddr0_wdata_i(41)
       , fabric_fpga_ddr0_wdata_i43                  =>  fabric_fpga_ddr0_wdata_i(42)
       , fabric_fpga_ddr0_wdata_i44                  =>  fabric_fpga_ddr0_wdata_i(43)
       , fabric_fpga_ddr0_wdata_i45                  =>  fabric_fpga_ddr0_wdata_i(44)
       , fabric_fpga_ddr0_wdata_i46                  =>  fabric_fpga_ddr0_wdata_i(45)
       , fabric_fpga_ddr0_wdata_i47                  =>  fabric_fpga_ddr0_wdata_i(46)
       , fabric_fpga_ddr0_wdata_i48                  =>  fabric_fpga_ddr0_wdata_i(47)
       , fabric_fpga_ddr0_wdata_i49                  =>  fabric_fpga_ddr0_wdata_i(48)
       , fabric_fpga_ddr0_wdata_i50                  =>  fabric_fpga_ddr0_wdata_i(49)
       , fabric_fpga_ddr0_wdata_i51                  =>  fabric_fpga_ddr0_wdata_i(50)
       , fabric_fpga_ddr0_wdata_i52                  =>  fabric_fpga_ddr0_wdata_i(51)
       , fabric_fpga_ddr0_wdata_i53                  =>  fabric_fpga_ddr0_wdata_i(52)
       , fabric_fpga_ddr0_wdata_i54                  =>  fabric_fpga_ddr0_wdata_i(53)
       , fabric_fpga_ddr0_wdata_i55                  =>  fabric_fpga_ddr0_wdata_i(54)
       , fabric_fpga_ddr0_wdata_i56                  =>  fabric_fpga_ddr0_wdata_i(55)
       , fabric_fpga_ddr0_wdata_i57                  =>  fabric_fpga_ddr0_wdata_i(56)
       , fabric_fpga_ddr0_wdata_i58                  =>  fabric_fpga_ddr0_wdata_i(57)
       , fabric_fpga_ddr0_wdata_i59                  =>  fabric_fpga_ddr0_wdata_i(58)
       , fabric_fpga_ddr0_wdata_i60                  =>  fabric_fpga_ddr0_wdata_i(59)
       , fabric_fpga_ddr0_wdata_i61                  =>  fabric_fpga_ddr0_wdata_i(60)
       , fabric_fpga_ddr0_wdata_i62                  =>  fabric_fpga_ddr0_wdata_i(61)
       , fabric_fpga_ddr0_wdata_i63                  =>  fabric_fpga_ddr0_wdata_i(62)
       , fabric_fpga_ddr0_wdata_i64                  =>  fabric_fpga_ddr0_wdata_i(63)
       , fabric_fpga_ddr0_wdata_i65                  =>  fabric_fpga_ddr0_wdata_i(64)
       , fabric_fpga_ddr0_wdata_i66                  =>  fabric_fpga_ddr0_wdata_i(65)
       , fabric_fpga_ddr0_wdata_i67                  =>  fabric_fpga_ddr0_wdata_i(66)
       , fabric_fpga_ddr0_wdata_i68                  =>  fabric_fpga_ddr0_wdata_i(67)
       , fabric_fpga_ddr0_wdata_i69                  =>  fabric_fpga_ddr0_wdata_i(68)
       , fabric_fpga_ddr0_wdata_i70                  =>  fabric_fpga_ddr0_wdata_i(69)
       , fabric_fpga_ddr0_wdata_i71                  =>  fabric_fpga_ddr0_wdata_i(70)
       , fabric_fpga_ddr0_wdata_i72                  =>  fabric_fpga_ddr0_wdata_i(71)
       , fabric_fpga_ddr0_wdata_i73                  =>  fabric_fpga_ddr0_wdata_i(72)
       , fabric_fpga_ddr0_wdata_i74                  =>  fabric_fpga_ddr0_wdata_i(73)
       , fabric_fpga_ddr0_wdata_i75                  =>  fabric_fpga_ddr0_wdata_i(74)
       , fabric_fpga_ddr0_wdata_i76                  =>  fabric_fpga_ddr0_wdata_i(75)
       , fabric_fpga_ddr0_wdata_i77                  =>  fabric_fpga_ddr0_wdata_i(76)
       , fabric_fpga_ddr0_wdata_i78                  =>  fabric_fpga_ddr0_wdata_i(77)
       , fabric_fpga_ddr0_wdata_i79                  =>  fabric_fpga_ddr0_wdata_i(78)
       , fabric_fpga_ddr0_wdata_i80                  =>  fabric_fpga_ddr0_wdata_i(79)
       , fabric_fpga_ddr0_wdata_i81                  =>  fabric_fpga_ddr0_wdata_i(80)
       , fabric_fpga_ddr0_wdata_i82                  =>  fabric_fpga_ddr0_wdata_i(81)
       , fabric_fpga_ddr0_wdata_i83                  =>  fabric_fpga_ddr0_wdata_i(82)
       , fabric_fpga_ddr0_wdata_i84                  =>  fabric_fpga_ddr0_wdata_i(83)
       , fabric_fpga_ddr0_wdata_i85                  =>  fabric_fpga_ddr0_wdata_i(84)
       , fabric_fpga_ddr0_wdata_i86                  =>  fabric_fpga_ddr0_wdata_i(85)
       , fabric_fpga_ddr0_wdata_i87                  =>  fabric_fpga_ddr0_wdata_i(86)
       , fabric_fpga_ddr0_wdata_i88                  =>  fabric_fpga_ddr0_wdata_i(87)
       , fabric_fpga_ddr0_wdata_i89                  =>  fabric_fpga_ddr0_wdata_i(88)
       , fabric_fpga_ddr0_wdata_i90                  =>  fabric_fpga_ddr0_wdata_i(89)
       , fabric_fpga_ddr0_wdata_i91                  =>  fabric_fpga_ddr0_wdata_i(90)
       , fabric_fpga_ddr0_wdata_i92                  =>  fabric_fpga_ddr0_wdata_i(91)
       , fabric_fpga_ddr0_wdata_i93                  =>  fabric_fpga_ddr0_wdata_i(92)
       , fabric_fpga_ddr0_wdata_i94                  =>  fabric_fpga_ddr0_wdata_i(93)
       , fabric_fpga_ddr0_wdata_i95                  =>  fabric_fpga_ddr0_wdata_i(94)
       , fabric_fpga_ddr0_wdata_i96                  =>  fabric_fpga_ddr0_wdata_i(95)
       , fabric_fpga_ddr0_wdata_i97                  =>  fabric_fpga_ddr0_wdata_i(96)
       , fabric_fpga_ddr0_wdata_i98                  =>  fabric_fpga_ddr0_wdata_i(97)
       , fabric_fpga_ddr0_wdata_i99                  =>  fabric_fpga_ddr0_wdata_i(98)
       , fabric_fpga_ddr0_wdata_i100                 =>  fabric_fpga_ddr0_wdata_i(99)
       , fabric_fpga_ddr0_wdata_i101                 =>  fabric_fpga_ddr0_wdata_i(100)
       , fabric_fpga_ddr0_wdata_i102                 =>  fabric_fpga_ddr0_wdata_i(101)
       , fabric_fpga_ddr0_wdata_i103                 =>  fabric_fpga_ddr0_wdata_i(102)
       , fabric_fpga_ddr0_wdata_i104                 =>  fabric_fpga_ddr0_wdata_i(103)
       , fabric_fpga_ddr0_wdata_i105                 =>  fabric_fpga_ddr0_wdata_i(104)
       , fabric_fpga_ddr0_wdata_i106                 =>  fabric_fpga_ddr0_wdata_i(105)
       , fabric_fpga_ddr0_wdata_i107                 =>  fabric_fpga_ddr0_wdata_i(106)
       , fabric_fpga_ddr0_wdata_i108                 =>  fabric_fpga_ddr0_wdata_i(107)
       , fabric_fpga_ddr0_wdata_i109                 =>  fabric_fpga_ddr0_wdata_i(108)
       , fabric_fpga_ddr0_wdata_i110                 =>  fabric_fpga_ddr0_wdata_i(109)
       , fabric_fpga_ddr0_wdata_i111                 =>  fabric_fpga_ddr0_wdata_i(110)
       , fabric_fpga_ddr0_wdata_i112                 =>  fabric_fpga_ddr0_wdata_i(111)
       , fabric_fpga_ddr0_wdata_i113                 =>  fabric_fpga_ddr0_wdata_i(112)
       , fabric_fpga_ddr0_wdata_i114                 =>  fabric_fpga_ddr0_wdata_i(113)
       , fabric_fpga_ddr0_wdata_i115                 =>  fabric_fpga_ddr0_wdata_i(114)
       , fabric_fpga_ddr0_wdata_i116                 =>  fabric_fpga_ddr0_wdata_i(115)
       , fabric_fpga_ddr0_wdata_i117                 =>  fabric_fpga_ddr0_wdata_i(116)
       , fabric_fpga_ddr0_wdata_i118                 =>  fabric_fpga_ddr0_wdata_i(117)
       , fabric_fpga_ddr0_wdata_i119                 =>  fabric_fpga_ddr0_wdata_i(118)
       , fabric_fpga_ddr0_wdata_i120                 =>  fabric_fpga_ddr0_wdata_i(119)
       , fabric_fpga_ddr0_wdata_i121                 =>  fabric_fpga_ddr0_wdata_i(120)
       , fabric_fpga_ddr0_wdata_i122                 =>  fabric_fpga_ddr0_wdata_i(121)
       , fabric_fpga_ddr0_wdata_i123                 =>  fabric_fpga_ddr0_wdata_i(122)
       , fabric_fpga_ddr0_wdata_i124                 =>  fabric_fpga_ddr0_wdata_i(123)
       , fabric_fpga_ddr0_wdata_i125                 =>  fabric_fpga_ddr0_wdata_i(124)
       , fabric_fpga_ddr0_wdata_i126                 =>  fabric_fpga_ddr0_wdata_i(125)
       , fabric_fpga_ddr0_wdata_i127                 =>  fabric_fpga_ddr0_wdata_i(126)
       , fabric_fpga_ddr0_wdata_i128                 =>  fabric_fpga_ddr0_wdata_i(127)
       , fabric_fpga_ddr0_wlast_i                    =>  fabric_fpga_ddr0_wlast_i
       , fabric_fpga_ddr0_wstrb_i1                   =>  fabric_fpga_ddr0_wstrb_i(0)
       , fabric_fpga_ddr0_wstrb_i2                   =>  fabric_fpga_ddr0_wstrb_i(1)
       , fabric_fpga_ddr0_wstrb_i3                   =>  fabric_fpga_ddr0_wstrb_i(2)
       , fabric_fpga_ddr0_wstrb_i4                   =>  fabric_fpga_ddr0_wstrb_i(3)
       , fabric_fpga_ddr0_wstrb_i5                   =>  fabric_fpga_ddr0_wstrb_i(4)
       , fabric_fpga_ddr0_wstrb_i6                   =>  fabric_fpga_ddr0_wstrb_i(5)
       , fabric_fpga_ddr0_wstrb_i7                   =>  fabric_fpga_ddr0_wstrb_i(6)
       , fabric_fpga_ddr0_wstrb_i8                   =>  fabric_fpga_ddr0_wstrb_i(7)
       , fabric_fpga_ddr0_wstrb_i9                   =>  fabric_fpga_ddr0_wstrb_i(8)
       , fabric_fpga_ddr0_wstrb_i10                  =>  fabric_fpga_ddr0_wstrb_i(9)
       , fabric_fpga_ddr0_wstrb_i11                  =>  fabric_fpga_ddr0_wstrb_i(10)
       , fabric_fpga_ddr0_wstrb_i12                  =>  fabric_fpga_ddr0_wstrb_i(11)
       , fabric_fpga_ddr0_wstrb_i13                  =>  fabric_fpga_ddr0_wstrb_i(12)
       , fabric_fpga_ddr0_wstrb_i14                  =>  fabric_fpga_ddr0_wstrb_i(13)
       , fabric_fpga_ddr0_wstrb_i15                  =>  fabric_fpga_ddr0_wstrb_i(14)
       , fabric_fpga_ddr0_wstrb_i16                  =>  fabric_fpga_ddr0_wstrb_i(15)
       , fabric_fpga_ddr0_wvalid_i                   =>  fabric_fpga_ddr0_wvalid_i
       , fabric_fpga_paddr_apb_o1                    =>  fabric_fpga_paddr_apb_o(0)
       , fabric_fpga_paddr_apb_o2                    =>  fabric_fpga_paddr_apb_o(1)
       , fabric_fpga_paddr_apb_o3                    =>  fabric_fpga_paddr_apb_o(2)
       , fabric_fpga_paddr_apb_o4                    =>  fabric_fpga_paddr_apb_o(3)
       , fabric_fpga_paddr_apb_o5                    =>  fabric_fpga_paddr_apb_o(4)
       , fabric_fpga_paddr_apb_o6                    =>  fabric_fpga_paddr_apb_o(5)
       , fabric_fpga_paddr_apb_o7                    =>  fabric_fpga_paddr_apb_o(6)
       , fabric_fpga_paddr_apb_o8                    =>  fabric_fpga_paddr_apb_o(7)
       , fabric_fpga_paddr_apb_o9                    =>  fabric_fpga_paddr_apb_o(8)
       , fabric_fpga_paddr_apb_o10                   =>  fabric_fpga_paddr_apb_o(9)
       , fabric_fpga_paddr_apb_o11                   =>  fabric_fpga_paddr_apb_o(10)
       , fabric_fpga_paddr_apb_o12                   =>  fabric_fpga_paddr_apb_o(11)
       , fabric_fpga_paddr_apb_o13                   =>  fabric_fpga_paddr_apb_o(12)
       , fabric_fpga_paddr_apb_o14                   =>  fabric_fpga_paddr_apb_o(13)
       , fabric_fpga_paddr_apb_o15                   =>  fabric_fpga_paddr_apb_o(14)
       , fabric_fpga_paddr_apb_o16                   =>  fabric_fpga_paddr_apb_o(15)
       , fabric_fpga_paddr_apb_o17                   =>  fabric_fpga_paddr_apb_o(16)
       , fabric_fpga_paddr_apb_o18                   =>  fabric_fpga_paddr_apb_o(17)
       , fabric_fpga_paddr_apb_o19                   =>  fabric_fpga_paddr_apb_o(18)
       , fabric_fpga_paddr_apb_o20                   =>  fabric_fpga_paddr_apb_o(19)
       , fabric_fpga_paddr_apb_o21                   =>  fabric_fpga_paddr_apb_o(20)
       , fabric_fpga_paddr_apb_o22                   =>  fabric_fpga_paddr_apb_o(21)
       , fabric_fpga_paddr_apb_o23                   =>  fabric_fpga_paddr_apb_o(22)
       , fabric_fpga_paddr_apb_o24                   =>  fabric_fpga_paddr_apb_o(23)
       , fabric_fpga_paddr_apb_o25                   =>  fabric_fpga_paddr_apb_o(24)
       , fabric_fpga_paddr_apb_o26                   =>  fabric_fpga_paddr_apb_o(25)
       , fabric_fpga_paddr_apb_o27                   =>  fabric_fpga_paddr_apb_o(26)
       , fabric_fpga_paddr_apb_o28                   =>  fabric_fpga_paddr_apb_o(27)
       , fabric_fpga_paddr_apb_o29                   =>  fabric_fpga_paddr_apb_o(28)
       , fabric_fpga_paddr_apb_o30                   =>  fabric_fpga_paddr_apb_o(29)
       , fabric_fpga_paddr_apb_o31                   =>  fabric_fpga_paddr_apb_o(30)
       , fabric_fpga_paddr_apb_o32                   =>  fabric_fpga_paddr_apb_o(31)
       , fabric_fpga_penable_apb_o                   =>  fabric_fpga_penable_apb_o
       , fabric_fpga_psel_apb_o                      =>  fabric_fpga_psel_apb_o
       , fabric_fpga_pwdata_apb_o1                   =>  fabric_fpga_pwdata_apb_o(0)
       , fabric_fpga_pwdata_apb_o2                   =>  fabric_fpga_pwdata_apb_o(1)
       , fabric_fpga_pwdata_apb_o3                   =>  fabric_fpga_pwdata_apb_o(2)
       , fabric_fpga_pwdata_apb_o4                   =>  fabric_fpga_pwdata_apb_o(3)
       , fabric_fpga_pwdata_apb_o5                   =>  fabric_fpga_pwdata_apb_o(4)
       , fabric_fpga_pwdata_apb_o6                   =>  fabric_fpga_pwdata_apb_o(5)
       , fabric_fpga_pwdata_apb_o7                   =>  fabric_fpga_pwdata_apb_o(6)
       , fabric_fpga_pwdata_apb_o8                   =>  fabric_fpga_pwdata_apb_o(7)
       , fabric_fpga_pwdata_apb_o9                   =>  fabric_fpga_pwdata_apb_o(8)
       , fabric_fpga_pwdata_apb_o10                  =>  fabric_fpga_pwdata_apb_o(9)
       , fabric_fpga_pwdata_apb_o11                  =>  fabric_fpga_pwdata_apb_o(10)
       , fabric_fpga_pwdata_apb_o12                  =>  fabric_fpga_pwdata_apb_o(11)
       , fabric_fpga_pwdata_apb_o13                  =>  fabric_fpga_pwdata_apb_o(12)
       , fabric_fpga_pwdata_apb_o14                  =>  fabric_fpga_pwdata_apb_o(13)
       , fabric_fpga_pwdata_apb_o15                  =>  fabric_fpga_pwdata_apb_o(14)
       , fabric_fpga_pwdata_apb_o16                  =>  fabric_fpga_pwdata_apb_o(15)
       , fabric_fpga_pwdata_apb_o17                  =>  fabric_fpga_pwdata_apb_o(16)
       , fabric_fpga_pwdata_apb_o18                  =>  fabric_fpga_pwdata_apb_o(17)
       , fabric_fpga_pwdata_apb_o19                  =>  fabric_fpga_pwdata_apb_o(18)
       , fabric_fpga_pwdata_apb_o20                  =>  fabric_fpga_pwdata_apb_o(19)
       , fabric_fpga_pwdata_apb_o21                  =>  fabric_fpga_pwdata_apb_o(20)
       , fabric_fpga_pwdata_apb_o22                  =>  fabric_fpga_pwdata_apb_o(21)
       , fabric_fpga_pwdata_apb_o23                  =>  fabric_fpga_pwdata_apb_o(22)
       , fabric_fpga_pwdata_apb_o24                  =>  fabric_fpga_pwdata_apb_o(23)
       , fabric_fpga_pwdata_apb_o25                  =>  fabric_fpga_pwdata_apb_o(24)
       , fabric_fpga_pwdata_apb_o26                  =>  fabric_fpga_pwdata_apb_o(25)
       , fabric_fpga_pwdata_apb_o27                  =>  fabric_fpga_pwdata_apb_o(26)
       , fabric_fpga_pwdata_apb_o28                  =>  fabric_fpga_pwdata_apb_o(27)
       , fabric_fpga_pwdata_apb_o29                  =>  fabric_fpga_pwdata_apb_o(28)
       , fabric_fpga_pwdata_apb_o30                  =>  fabric_fpga_pwdata_apb_o(29)
       , fabric_fpga_pwdata_apb_o31                  =>  fabric_fpga_pwdata_apb_o(30)
       , fabric_fpga_pwdata_apb_o32                  =>  fabric_fpga_pwdata_apb_o(31)
       , fabric_fpga_pwrite_apb_o                    =>  fabric_fpga_pwrite_apb_o
       , fabric_fpga_prdata_apb_i1                   =>  fabric_fpga_prdata_apb_i(0)
       , fabric_fpga_prdata_apb_i2                   =>  fabric_fpga_prdata_apb_i(1)
       , fabric_fpga_prdata_apb_i3                   =>  fabric_fpga_prdata_apb_i(2)
       , fabric_fpga_prdata_apb_i4                   =>  fabric_fpga_prdata_apb_i(3)
       , fabric_fpga_prdata_apb_i5                   =>  fabric_fpga_prdata_apb_i(4)
       , fabric_fpga_prdata_apb_i6                   =>  fabric_fpga_prdata_apb_i(5)
       , fabric_fpga_prdata_apb_i7                   =>  fabric_fpga_prdata_apb_i(6)
       , fabric_fpga_prdata_apb_i8                   =>  fabric_fpga_prdata_apb_i(7)
       , fabric_fpga_prdata_apb_i9                   =>  fabric_fpga_prdata_apb_i(8)
       , fabric_fpga_prdata_apb_i10                  =>  fabric_fpga_prdata_apb_i(9)
       , fabric_fpga_prdata_apb_i11                  =>  fabric_fpga_prdata_apb_i(10)
       , fabric_fpga_prdata_apb_i12                  =>  fabric_fpga_prdata_apb_i(11)
       , fabric_fpga_prdata_apb_i13                  =>  fabric_fpga_prdata_apb_i(12)
       , fabric_fpga_prdata_apb_i14                  =>  fabric_fpga_prdata_apb_i(13)
       , fabric_fpga_prdata_apb_i15                  =>  fabric_fpga_prdata_apb_i(14)
       , fabric_fpga_prdata_apb_i16                  =>  fabric_fpga_prdata_apb_i(15)
       , fabric_fpga_prdata_apb_i17                  =>  fabric_fpga_prdata_apb_i(16)
       , fabric_fpga_prdata_apb_i18                  =>  fabric_fpga_prdata_apb_i(17)
       , fabric_fpga_prdata_apb_i19                  =>  fabric_fpga_prdata_apb_i(18)
       , fabric_fpga_prdata_apb_i20                  =>  fabric_fpga_prdata_apb_i(19)
       , fabric_fpga_prdata_apb_i21                  =>  fabric_fpga_prdata_apb_i(20)
       , fabric_fpga_prdata_apb_i22                  =>  fabric_fpga_prdata_apb_i(21)
       , fabric_fpga_prdata_apb_i23                  =>  fabric_fpga_prdata_apb_i(22)
       , fabric_fpga_prdata_apb_i24                  =>  fabric_fpga_prdata_apb_i(23)
       , fabric_fpga_prdata_apb_i25                  =>  fabric_fpga_prdata_apb_i(24)
       , fabric_fpga_prdata_apb_i26                  =>  fabric_fpga_prdata_apb_i(25)
       , fabric_fpga_prdata_apb_i27                  =>  fabric_fpga_prdata_apb_i(26)
       , fabric_fpga_prdata_apb_i28                  =>  fabric_fpga_prdata_apb_i(27)
       , fabric_fpga_prdata_apb_i29                  =>  fabric_fpga_prdata_apb_i(28)
       , fabric_fpga_prdata_apb_i30                  =>  fabric_fpga_prdata_apb_i(29)
       , fabric_fpga_prdata_apb_i31                  =>  fabric_fpga_prdata_apb_i(30)
       , fabric_fpga_prdata_apb_i32                  =>  fabric_fpga_prdata_apb_i(31)
       , fabric_fpga_pready_apb_i                    =>  fabric_fpga_pready_apb_i
       , fabric_fpga_pslverr_apb_i                   =>  fabric_fpga_pslverr_apb_i
       , fabric_llpp0_araddr_s_o1                    =>  fabric_llpp0_araddr_s_o(0)
       , fabric_llpp0_araddr_s_o2                    =>  fabric_llpp0_araddr_s_o(1)
       , fabric_llpp0_araddr_s_o3                    =>  fabric_llpp0_araddr_s_o(2)
       , fabric_llpp0_araddr_s_o4                    =>  fabric_llpp0_araddr_s_o(3)
       , fabric_llpp0_araddr_s_o5                    =>  fabric_llpp0_araddr_s_o(4)
       , fabric_llpp0_araddr_s_o6                    =>  fabric_llpp0_araddr_s_o(5)
       , fabric_llpp0_araddr_s_o7                    =>  fabric_llpp0_araddr_s_o(6)
       , fabric_llpp0_araddr_s_o8                    =>  fabric_llpp0_araddr_s_o(7)
       , fabric_llpp0_araddr_s_o9                    =>  fabric_llpp0_araddr_s_o(8)
       , fabric_llpp0_araddr_s_o10                   =>  fabric_llpp0_araddr_s_o(9)
       , fabric_llpp0_araddr_s_o11                   =>  fabric_llpp0_araddr_s_o(10)
       , fabric_llpp0_araddr_s_o12                   =>  fabric_llpp0_araddr_s_o(11)
       , fabric_llpp0_araddr_s_o13                   =>  fabric_llpp0_araddr_s_o(12)
       , fabric_llpp0_araddr_s_o14                   =>  fabric_llpp0_araddr_s_o(13)
       , fabric_llpp0_araddr_s_o15                   =>  fabric_llpp0_araddr_s_o(14)
       , fabric_llpp0_araddr_s_o16                   =>  fabric_llpp0_araddr_s_o(15)
       , fabric_llpp0_araddr_s_o17                   =>  fabric_llpp0_araddr_s_o(16)
       , fabric_llpp0_araddr_s_o18                   =>  fabric_llpp0_araddr_s_o(17)
       , fabric_llpp0_araddr_s_o19                   =>  fabric_llpp0_araddr_s_o(18)
       , fabric_llpp0_araddr_s_o20                   =>  fabric_llpp0_araddr_s_o(19)
       , fabric_llpp0_araddr_s_o21                   =>  fabric_llpp0_araddr_s_o(20)
       , fabric_llpp0_araddr_s_o22                   =>  fabric_llpp0_araddr_s_o(21)
       , fabric_llpp0_araddr_s_o23                   =>  fabric_llpp0_araddr_s_o(22)
       , fabric_llpp0_araddr_s_o24                   =>  fabric_llpp0_araddr_s_o(23)
       , fabric_llpp0_araddr_s_o25                   =>  fabric_llpp0_araddr_s_o(24)
       , fabric_llpp0_araddr_s_o26                   =>  fabric_llpp0_araddr_s_o(25)
       , fabric_llpp0_araddr_s_o27                   =>  fabric_llpp0_araddr_s_o(26)
       , fabric_llpp0_araddr_s_o28                   =>  fabric_llpp0_araddr_s_o(27)
       , fabric_llpp0_araddr_s_o29                   =>  fabric_llpp0_araddr_s_o(28)
       , fabric_llpp0_araddr_s_o30                   =>  fabric_llpp0_araddr_s_o(29)
       , fabric_llpp0_araddr_s_o31                   =>  fabric_llpp0_araddr_s_o(30)
       , fabric_llpp0_araddr_s_o32                   =>  fabric_llpp0_araddr_s_o(31)
       , fabric_llpp0_arburst_s_o1                   =>  fabric_llpp0_arburst_s_o(0)
       , fabric_llpp0_arburst_s_o2                   =>  fabric_llpp0_arburst_s_o(1)
       , fabric_llpp0_arcache_s_o1                   =>  fabric_llpp0_arcache_s_o(0)
       , fabric_llpp0_arcache_s_o2                   =>  fabric_llpp0_arcache_s_o(1)
       , fabric_llpp0_arcache_s_o3                   =>  fabric_llpp0_arcache_s_o(2)
       , fabric_llpp0_arcache_s_o4                   =>  fabric_llpp0_arcache_s_o(3)
       , fabric_llpp0_arid_s_o1                      =>  fabric_llpp0_arid_s_o(0)
       , fabric_llpp0_arid_s_o2                      =>  fabric_llpp0_arid_s_o(1)
       , fabric_llpp0_arid_s_o3                      =>  fabric_llpp0_arid_s_o(2)
       , fabric_llpp0_arid_s_o4                      =>  fabric_llpp0_arid_s_o(3)
       , fabric_llpp0_arid_s_o5                      =>  fabric_llpp0_arid_s_o(4)
       , fabric_llpp0_arid_s_o6                      =>  fabric_llpp0_arid_s_o(5)
       , fabric_llpp0_arid_s_o7                      =>  fabric_llpp0_arid_s_o(6)
       , fabric_llpp0_arid_s_o8                      =>  fabric_llpp0_arid_s_o(7)
       , fabric_llpp0_arid_s_o9                      =>  fabric_llpp0_arid_s_o(8)
       , fabric_llpp0_arid_s_o10                     =>  fabric_llpp0_arid_s_o(9)
       , fabric_llpp0_arid_s_o11                     =>  fabric_llpp0_arid_s_o(10)
       , fabric_llpp0_arid_s_o12                     =>  fabric_llpp0_arid_s_o(11)
       , fabric_llpp0_arlen_s_o1                     =>  fabric_llpp0_arlen_s_o(0)
       , fabric_llpp0_arlen_s_o2                     =>  fabric_llpp0_arlen_s_o(1)
       , fabric_llpp0_arlen_s_o3                     =>  fabric_llpp0_arlen_s_o(2)
       , fabric_llpp0_arlen_s_o4                     =>  fabric_llpp0_arlen_s_o(3)
       , fabric_llpp0_arlen_s_o5                     =>  fabric_llpp0_arlen_s_o(4)
       , fabric_llpp0_arlen_s_o6                     =>  fabric_llpp0_arlen_s_o(5)
       , fabric_llpp0_arlen_s_o7                     =>  fabric_llpp0_arlen_s_o(6)
       , fabric_llpp0_arlen_s_o8                     =>  fabric_llpp0_arlen_s_o(7)
       , fabric_llpp0_arlock_s_o                     =>  fabric_llpp0_arlock_s_o
       , fabric_llpp0_arprot_s_o1                    =>  fabric_llpp0_arprot_s_o(0)
       , fabric_llpp0_arprot_s_o2                    =>  fabric_llpp0_arprot_s_o(1)
       , fabric_llpp0_arprot_s_o3                    =>  fabric_llpp0_arprot_s_o(2)
       , fabric_llpp0_arqos_s_o1                     =>  fabric_llpp0_arqos_s_o(0)
       , fabric_llpp0_arqos_s_o2                     =>  fabric_llpp0_arqos_s_o(1)
       , fabric_llpp0_arqos_s_o3                     =>  fabric_llpp0_arqos_s_o(2)
       , fabric_llpp0_arqos_s_o4                     =>  fabric_llpp0_arqos_s_o(3)
       , fabric_llpp0_arsize_s_o1                    =>  fabric_llpp0_arsize_s_o(0)
       , fabric_llpp0_arsize_s_o2                    =>  fabric_llpp0_arsize_s_o(1)
       , fabric_llpp0_arsize_s_o3                    =>  fabric_llpp0_arsize_s_o(2)
       , fabric_llpp0_arvalid_s_o                    =>  fabric_llpp0_arvalid_s_o
       , fabric_llpp0_awaddr_s_o1                    =>  fabric_llpp0_awaddr_s_o(0)
       , fabric_llpp0_awaddr_s_o2                    =>  fabric_llpp0_awaddr_s_o(1)
       , fabric_llpp0_awaddr_s_o3                    =>  fabric_llpp0_awaddr_s_o(2)
       , fabric_llpp0_awaddr_s_o4                    =>  fabric_llpp0_awaddr_s_o(3)
       , fabric_llpp0_awaddr_s_o5                    =>  fabric_llpp0_awaddr_s_o(4)
       , fabric_llpp0_awaddr_s_o6                    =>  fabric_llpp0_awaddr_s_o(5)
       , fabric_llpp0_awaddr_s_o7                    =>  fabric_llpp0_awaddr_s_o(6)
       , fabric_llpp0_awaddr_s_o8                    =>  fabric_llpp0_awaddr_s_o(7)
       , fabric_llpp0_awaddr_s_o9                    =>  fabric_llpp0_awaddr_s_o(8)
       , fabric_llpp0_awaddr_s_o10                   =>  fabric_llpp0_awaddr_s_o(9)
       , fabric_llpp0_awaddr_s_o11                   =>  fabric_llpp0_awaddr_s_o(10)
       , fabric_llpp0_awaddr_s_o12                   =>  fabric_llpp0_awaddr_s_o(11)
       , fabric_llpp0_awaddr_s_o13                   =>  fabric_llpp0_awaddr_s_o(12)
       , fabric_llpp0_awaddr_s_o14                   =>  fabric_llpp0_awaddr_s_o(13)
       , fabric_llpp0_awaddr_s_o15                   =>  fabric_llpp0_awaddr_s_o(14)
       , fabric_llpp0_awaddr_s_o16                   =>  fabric_llpp0_awaddr_s_o(15)
       , fabric_llpp0_awaddr_s_o17                   =>  fabric_llpp0_awaddr_s_o(16)
       , fabric_llpp0_awaddr_s_o18                   =>  fabric_llpp0_awaddr_s_o(17)
       , fabric_llpp0_awaddr_s_o19                   =>  fabric_llpp0_awaddr_s_o(18)
       , fabric_llpp0_awaddr_s_o20                   =>  fabric_llpp0_awaddr_s_o(19)
       , fabric_llpp0_awaddr_s_o21                   =>  fabric_llpp0_awaddr_s_o(20)
       , fabric_llpp0_awaddr_s_o22                   =>  fabric_llpp0_awaddr_s_o(21)
       , fabric_llpp0_awaddr_s_o23                   =>  fabric_llpp0_awaddr_s_o(22)
       , fabric_llpp0_awaddr_s_o24                   =>  fabric_llpp0_awaddr_s_o(23)
       , fabric_llpp0_awaddr_s_o25                   =>  fabric_llpp0_awaddr_s_o(24)
       , fabric_llpp0_awaddr_s_o26                   =>  fabric_llpp0_awaddr_s_o(25)
       , fabric_llpp0_awaddr_s_o27                   =>  fabric_llpp0_awaddr_s_o(26)
       , fabric_llpp0_awaddr_s_o28                   =>  fabric_llpp0_awaddr_s_o(27)
       , fabric_llpp0_awaddr_s_o29                   =>  fabric_llpp0_awaddr_s_o(28)
       , fabric_llpp0_awaddr_s_o30                   =>  fabric_llpp0_awaddr_s_o(29)
       , fabric_llpp0_awaddr_s_o31                   =>  fabric_llpp0_awaddr_s_o(30)
       , fabric_llpp0_awaddr_s_o32                   =>  fabric_llpp0_awaddr_s_o(31)
       , fabric_llpp0_awburst_s_o1                   =>  fabric_llpp0_awburst_s_o(0)
       , fabric_llpp0_awburst_s_o2                   =>  fabric_llpp0_awburst_s_o(1)
       , fabric_llpp0_awcache_s_o1                   =>  fabric_llpp0_awcache_s_o(0)
       , fabric_llpp0_awcache_s_o2                   =>  fabric_llpp0_awcache_s_o(1)
       , fabric_llpp0_awcache_s_o3                   =>  fabric_llpp0_awcache_s_o(2)
       , fabric_llpp0_awcache_s_o4                   =>  fabric_llpp0_awcache_s_o(3)
       , fabric_llpp0_awid_s_o1                      =>  fabric_llpp0_awid_s_o(0)
       , fabric_llpp0_awid_s_o2                      =>  fabric_llpp0_awid_s_o(1)
       , fabric_llpp0_awid_s_o3                      =>  fabric_llpp0_awid_s_o(2)
       , fabric_llpp0_awid_s_o4                      =>  fabric_llpp0_awid_s_o(3)
       , fabric_llpp0_awid_s_o5                      =>  fabric_llpp0_awid_s_o(4)
       , fabric_llpp0_awid_s_o6                      =>  fabric_llpp0_awid_s_o(5)
       , fabric_llpp0_awid_s_o7                      =>  fabric_llpp0_awid_s_o(6)
       , fabric_llpp0_awid_s_o8                      =>  fabric_llpp0_awid_s_o(7)
       , fabric_llpp0_awid_s_o9                      =>  fabric_llpp0_awid_s_o(8)
       , fabric_llpp0_awid_s_o10                     =>  fabric_llpp0_awid_s_o(9)
       , fabric_llpp0_awid_s_o11                     =>  fabric_llpp0_awid_s_o(10)
       , fabric_llpp0_awid_s_o12                     =>  fabric_llpp0_awid_s_o(11)
       , fabric_llpp0_awlen_s_o1                     =>  fabric_llpp0_awlen_s_o(0)
       , fabric_llpp0_awlen_s_o2                     =>  fabric_llpp0_awlen_s_o(1)
       , fabric_llpp0_awlen_s_o3                     =>  fabric_llpp0_awlen_s_o(2)
       , fabric_llpp0_awlen_s_o4                     =>  fabric_llpp0_awlen_s_o(3)
       , fabric_llpp0_awlen_s_o5                     =>  fabric_llpp0_awlen_s_o(4)
       , fabric_llpp0_awlen_s_o6                     =>  fabric_llpp0_awlen_s_o(5)
       , fabric_llpp0_awlen_s_o7                     =>  fabric_llpp0_awlen_s_o(6)
       , fabric_llpp0_awlen_s_o8                     =>  fabric_llpp0_awlen_s_o(7)
       , fabric_llpp0_awlock_s_o                     =>  fabric_llpp0_awlock_s_o
       , fabric_llpp0_awprot_s_o1                    =>  fabric_llpp0_awprot_s_o(0)
       , fabric_llpp0_awprot_s_o2                    =>  fabric_llpp0_awprot_s_o(1)
       , fabric_llpp0_awprot_s_o3                    =>  fabric_llpp0_awprot_s_o(2)
       , fabric_llpp0_awqos_s_o1                     =>  fabric_llpp0_awqos_s_o(0)
       , fabric_llpp0_awqos_s_o2                     =>  fabric_llpp0_awqos_s_o(1)
       , fabric_llpp0_awqos_s_o3                     =>  fabric_llpp0_awqos_s_o(2)
       , fabric_llpp0_awqos_s_o4                     =>  fabric_llpp0_awqos_s_o(3)
       , fabric_llpp0_awsize_s_o1                    =>  fabric_llpp0_awsize_s_o(0)
       , fabric_llpp0_awsize_s_o2                    =>  fabric_llpp0_awsize_s_o(1)
       , fabric_llpp0_awsize_s_o3                    =>  fabric_llpp0_awsize_s_o(2)
       , fabric_llpp0_awvalid_s_o                    =>  fabric_llpp0_awvalid_s_o
       , fabric_llpp0_bready_s_o                     =>  fabric_llpp0_bready_s_o
       , fabric_llpp0_rready_s_o                     =>  fabric_llpp0_rready_s_o
       , fabric_llpp0_wdata_s_o1                     =>  fabric_llpp0_wdata_s_o(0)
       , fabric_llpp0_wdata_s_o2                     =>  fabric_llpp0_wdata_s_o(1)
       , fabric_llpp0_wdata_s_o3                     =>  fabric_llpp0_wdata_s_o(2)
       , fabric_llpp0_wdata_s_o4                     =>  fabric_llpp0_wdata_s_o(3)
       , fabric_llpp0_wdata_s_o5                     =>  fabric_llpp0_wdata_s_o(4)
       , fabric_llpp0_wdata_s_o6                     =>  fabric_llpp0_wdata_s_o(5)
       , fabric_llpp0_wdata_s_o7                     =>  fabric_llpp0_wdata_s_o(6)
       , fabric_llpp0_wdata_s_o8                     =>  fabric_llpp0_wdata_s_o(7)
       , fabric_llpp0_wdata_s_o9                     =>  fabric_llpp0_wdata_s_o(8)
       , fabric_llpp0_wdata_s_o10                    =>  fabric_llpp0_wdata_s_o(9)
       , fabric_llpp0_wdata_s_o11                    =>  fabric_llpp0_wdata_s_o(10)
       , fabric_llpp0_wdata_s_o12                    =>  fabric_llpp0_wdata_s_o(11)
       , fabric_llpp0_wdata_s_o13                    =>  fabric_llpp0_wdata_s_o(12)
       , fabric_llpp0_wdata_s_o14                    =>  fabric_llpp0_wdata_s_o(13)
       , fabric_llpp0_wdata_s_o15                    =>  fabric_llpp0_wdata_s_o(14)
       , fabric_llpp0_wdata_s_o16                    =>  fabric_llpp0_wdata_s_o(15)
       , fabric_llpp0_wdata_s_o17                    =>  fabric_llpp0_wdata_s_o(16)
       , fabric_llpp0_wdata_s_o18                    =>  fabric_llpp0_wdata_s_o(17)
       , fabric_llpp0_wdata_s_o19                    =>  fabric_llpp0_wdata_s_o(18)
       , fabric_llpp0_wdata_s_o20                    =>  fabric_llpp0_wdata_s_o(19)
       , fabric_llpp0_wdata_s_o21                    =>  fabric_llpp0_wdata_s_o(20)
       , fabric_llpp0_wdata_s_o22                    =>  fabric_llpp0_wdata_s_o(21)
       , fabric_llpp0_wdata_s_o23                    =>  fabric_llpp0_wdata_s_o(22)
       , fabric_llpp0_wdata_s_o24                    =>  fabric_llpp0_wdata_s_o(23)
       , fabric_llpp0_wdata_s_o25                    =>  fabric_llpp0_wdata_s_o(24)
       , fabric_llpp0_wdata_s_o26                    =>  fabric_llpp0_wdata_s_o(25)
       , fabric_llpp0_wdata_s_o27                    =>  fabric_llpp0_wdata_s_o(26)
       , fabric_llpp0_wdata_s_o28                    =>  fabric_llpp0_wdata_s_o(27)
       , fabric_llpp0_wdata_s_o29                    =>  fabric_llpp0_wdata_s_o(28)
       , fabric_llpp0_wdata_s_o30                    =>  fabric_llpp0_wdata_s_o(29)
       , fabric_llpp0_wdata_s_o31                    =>  fabric_llpp0_wdata_s_o(30)
       , fabric_llpp0_wdata_s_o32                    =>  fabric_llpp0_wdata_s_o(31)
       , fabric_llpp0_wlast_s_o                      =>  fabric_llpp0_wlast_s_o
       , fabric_llpp0_wstrb_s_o1                     =>  fabric_llpp0_wstrb_s_o(0)
       , fabric_llpp0_wstrb_s_o2                     =>  fabric_llpp0_wstrb_s_o(1)
       , fabric_llpp0_wstrb_s_o3                     =>  fabric_llpp0_wstrb_s_o(2)
       , fabric_llpp0_wstrb_s_o4                     =>  fabric_llpp0_wstrb_s_o(3)
       , fabric_llpp0_wvalid_s_o                     =>  fabric_llpp0_wvalid_s_o
       , fabric_llpp0_arready_s_i                    =>  fabric_llpp0_arready_s_i
       , fabric_llpp0_awready_s_i                    =>  fabric_llpp0_awready_s_i
       , fabric_llpp0_bid_s_i1                       =>  fabric_llpp0_bid_s_i(0)
       , fabric_llpp0_bid_s_i2                       =>  fabric_llpp0_bid_s_i(1)
       , fabric_llpp0_bid_s_i3                       =>  fabric_llpp0_bid_s_i(2)
       , fabric_llpp0_bid_s_i4                       =>  fabric_llpp0_bid_s_i(3)
       , fabric_llpp0_bid_s_i5                       =>  fabric_llpp0_bid_s_i(4)
       , fabric_llpp0_bid_s_i6                       =>  fabric_llpp0_bid_s_i(5)
       , fabric_llpp0_bid_s_i7                       =>  fabric_llpp0_bid_s_i(6)
       , fabric_llpp0_bid_s_i8                       =>  fabric_llpp0_bid_s_i(7)
       , fabric_llpp0_bid_s_i9                       =>  fabric_llpp0_bid_s_i(8)
       , fabric_llpp0_bid_s_i10                      =>  fabric_llpp0_bid_s_i(9)
       , fabric_llpp0_bid_s_i11                      =>  fabric_llpp0_bid_s_i(10)
       , fabric_llpp0_bid_s_i12                      =>  fabric_llpp0_bid_s_i(11)
       , fabric_llpp0_bresp_s_i1                     =>  fabric_llpp0_bresp_s_i(0)
       , fabric_llpp0_bresp_s_i2                     =>  fabric_llpp0_bresp_s_i(1)
       , fabric_llpp0_bvalid_s_i                     =>  fabric_llpp0_bvalid_s_i
       , fabric_llpp0_rdata_s_i1                     =>  fabric_llpp0_rdata_s_i(0)
       , fabric_llpp0_rdata_s_i2                     =>  fabric_llpp0_rdata_s_i(1)
       , fabric_llpp0_rdata_s_i3                     =>  fabric_llpp0_rdata_s_i(2)
       , fabric_llpp0_rdata_s_i4                     =>  fabric_llpp0_rdata_s_i(3)
       , fabric_llpp0_rdata_s_i5                     =>  fabric_llpp0_rdata_s_i(4)
       , fabric_llpp0_rdata_s_i6                     =>  fabric_llpp0_rdata_s_i(5)
       , fabric_llpp0_rdata_s_i7                     =>  fabric_llpp0_rdata_s_i(6)
       , fabric_llpp0_rdata_s_i8                     =>  fabric_llpp0_rdata_s_i(7)
       , fabric_llpp0_rdata_s_i9                     =>  fabric_llpp0_rdata_s_i(8)
       , fabric_llpp0_rdata_s_i10                    =>  fabric_llpp0_rdata_s_i(9)
       , fabric_llpp0_rdata_s_i11                    =>  fabric_llpp0_rdata_s_i(10)
       , fabric_llpp0_rdata_s_i12                    =>  fabric_llpp0_rdata_s_i(11)
       , fabric_llpp0_rdata_s_i13                    =>  fabric_llpp0_rdata_s_i(12)
       , fabric_llpp0_rdata_s_i14                    =>  fabric_llpp0_rdata_s_i(13)
       , fabric_llpp0_rdata_s_i15                    =>  fabric_llpp0_rdata_s_i(14)
       , fabric_llpp0_rdata_s_i16                    =>  fabric_llpp0_rdata_s_i(15)
       , fabric_llpp0_rdata_s_i17                    =>  fabric_llpp0_rdata_s_i(16)
       , fabric_llpp0_rdata_s_i18                    =>  fabric_llpp0_rdata_s_i(17)
       , fabric_llpp0_rdata_s_i19                    =>  fabric_llpp0_rdata_s_i(18)
       , fabric_llpp0_rdata_s_i20                    =>  fabric_llpp0_rdata_s_i(19)
       , fabric_llpp0_rdata_s_i21                    =>  fabric_llpp0_rdata_s_i(20)
       , fabric_llpp0_rdata_s_i22                    =>  fabric_llpp0_rdata_s_i(21)
       , fabric_llpp0_rdata_s_i23                    =>  fabric_llpp0_rdata_s_i(22)
       , fabric_llpp0_rdata_s_i24                    =>  fabric_llpp0_rdata_s_i(23)
       , fabric_llpp0_rdata_s_i25                    =>  fabric_llpp0_rdata_s_i(24)
       , fabric_llpp0_rdata_s_i26                    =>  fabric_llpp0_rdata_s_i(25)
       , fabric_llpp0_rdata_s_i27                    =>  fabric_llpp0_rdata_s_i(26)
       , fabric_llpp0_rdata_s_i28                    =>  fabric_llpp0_rdata_s_i(27)
       , fabric_llpp0_rdata_s_i29                    =>  fabric_llpp0_rdata_s_i(28)
       , fabric_llpp0_rdata_s_i30                    =>  fabric_llpp0_rdata_s_i(29)
       , fabric_llpp0_rdata_s_i31                    =>  fabric_llpp0_rdata_s_i(30)
       , fabric_llpp0_rdata_s_i32                    =>  fabric_llpp0_rdata_s_i(31)
       , fabric_llpp0_rid_s_i1                       =>  fabric_llpp0_rid_s_i(0)
       , fabric_llpp0_rid_s_i2                       =>  fabric_llpp0_rid_s_i(1)
       , fabric_llpp0_rid_s_i3                       =>  fabric_llpp0_rid_s_i(2)
       , fabric_llpp0_rid_s_i4                       =>  fabric_llpp0_rid_s_i(3)
       , fabric_llpp0_rid_s_i5                       =>  fabric_llpp0_rid_s_i(4)
       , fabric_llpp0_rid_s_i6                       =>  fabric_llpp0_rid_s_i(5)
       , fabric_llpp0_rid_s_i7                       =>  fabric_llpp0_rid_s_i(6)
       , fabric_llpp0_rid_s_i8                       =>  fabric_llpp0_rid_s_i(7)
       , fabric_llpp0_rid_s_i9                       =>  fabric_llpp0_rid_s_i(8)
       , fabric_llpp0_rid_s_i10                      =>  fabric_llpp0_rid_s_i(9)
       , fabric_llpp0_rid_s_i11                      =>  fabric_llpp0_rid_s_i(10)
       , fabric_llpp0_rid_s_i12                      =>  fabric_llpp0_rid_s_i(11)
       , fabric_llpp0_rlast_s_i                      =>  fabric_llpp0_rlast_s_i
       , fabric_llpp0_rresp_s_i1                     =>  fabric_llpp0_rresp_s_i(0)
       , fabric_llpp0_rresp_s_i2                     =>  fabric_llpp0_rresp_s_i(1)
       , fabric_llpp0_rvalid_s_i                     =>  fabric_llpp0_rvalid_s_i
       , fabric_llpp0_wready_s_i                     =>  fabric_llpp0_wready_s_i
       , fabric_llpp1_araddr_s_o1                    =>  fabric_llpp1_araddr_s_o(0)
       , fabric_llpp1_araddr_s_o2                    =>  fabric_llpp1_araddr_s_o(1)
       , fabric_llpp1_araddr_s_o3                    =>  fabric_llpp1_araddr_s_o(2)
       , fabric_llpp1_araddr_s_o4                    =>  fabric_llpp1_araddr_s_o(3)
       , fabric_llpp1_araddr_s_o5                    =>  fabric_llpp1_araddr_s_o(4)
       , fabric_llpp1_araddr_s_o6                    =>  fabric_llpp1_araddr_s_o(5)
       , fabric_llpp1_araddr_s_o7                    =>  fabric_llpp1_araddr_s_o(6)
       , fabric_llpp1_araddr_s_o8                    =>  fabric_llpp1_araddr_s_o(7)
       , fabric_llpp1_araddr_s_o9                    =>  fabric_llpp1_araddr_s_o(8)
       , fabric_llpp1_araddr_s_o10                   =>  fabric_llpp1_araddr_s_o(9)
       , fabric_llpp1_araddr_s_o11                   =>  fabric_llpp1_araddr_s_o(10)
       , fabric_llpp1_araddr_s_o12                   =>  fabric_llpp1_araddr_s_o(11)
       , fabric_llpp1_araddr_s_o13                   =>  fabric_llpp1_araddr_s_o(12)
       , fabric_llpp1_araddr_s_o14                   =>  fabric_llpp1_araddr_s_o(13)
       , fabric_llpp1_araddr_s_o15                   =>  fabric_llpp1_araddr_s_o(14)
       , fabric_llpp1_araddr_s_o16                   =>  fabric_llpp1_araddr_s_o(15)
       , fabric_llpp1_araddr_s_o17                   =>  fabric_llpp1_araddr_s_o(16)
       , fabric_llpp1_araddr_s_o18                   =>  fabric_llpp1_araddr_s_o(17)
       , fabric_llpp1_araddr_s_o19                   =>  fabric_llpp1_araddr_s_o(18)
       , fabric_llpp1_araddr_s_o20                   =>  fabric_llpp1_araddr_s_o(19)
       , fabric_llpp1_araddr_s_o21                   =>  fabric_llpp1_araddr_s_o(20)
       , fabric_llpp1_araddr_s_o22                   =>  fabric_llpp1_araddr_s_o(21)
       , fabric_llpp1_araddr_s_o23                   =>  fabric_llpp1_araddr_s_o(22)
       , fabric_llpp1_araddr_s_o24                   =>  fabric_llpp1_araddr_s_o(23)
       , fabric_llpp1_araddr_s_o25                   =>  fabric_llpp1_araddr_s_o(24)
       , fabric_llpp1_araddr_s_o26                   =>  fabric_llpp1_araddr_s_o(25)
       , fabric_llpp1_araddr_s_o27                   =>  fabric_llpp1_araddr_s_o(26)
       , fabric_llpp1_araddr_s_o28                   =>  fabric_llpp1_araddr_s_o(27)
       , fabric_llpp1_araddr_s_o29                   =>  fabric_llpp1_araddr_s_o(28)
       , fabric_llpp1_araddr_s_o30                   =>  fabric_llpp1_araddr_s_o(29)
       , fabric_llpp1_araddr_s_o31                   =>  fabric_llpp1_araddr_s_o(30)
       , fabric_llpp1_araddr_s_o32                   =>  fabric_llpp1_araddr_s_o(31)
       , fabric_llpp1_arburst_s_o1                   =>  fabric_llpp1_arburst_s_o(0)
       , fabric_llpp1_arburst_s_o2                   =>  fabric_llpp1_arburst_s_o(1)
       , fabric_llpp1_arcache_s_o1                   =>  fabric_llpp1_arcache_s_o(0)
       , fabric_llpp1_arcache_s_o2                   =>  fabric_llpp1_arcache_s_o(1)
       , fabric_llpp1_arcache_s_o3                   =>  fabric_llpp1_arcache_s_o(2)
       , fabric_llpp1_arcache_s_o4                   =>  fabric_llpp1_arcache_s_o(3)
       , fabric_llpp1_arid_s_o1                      =>  fabric_llpp1_arid_s_o(0)
       , fabric_llpp1_arid_s_o2                      =>  fabric_llpp1_arid_s_o(1)
       , fabric_llpp1_arid_s_o3                      =>  fabric_llpp1_arid_s_o(2)
       , fabric_llpp1_arid_s_o4                      =>  fabric_llpp1_arid_s_o(3)
       , fabric_llpp1_arid_s_o5                      =>  fabric_llpp1_arid_s_o(4)
       , fabric_llpp1_arid_s_o6                      =>  fabric_llpp1_arid_s_o(5)
       , fabric_llpp1_arid_s_o7                      =>  fabric_llpp1_arid_s_o(6)
       , fabric_llpp1_arid_s_o8                      =>  fabric_llpp1_arid_s_o(7)
       , fabric_llpp1_arid_s_o9                      =>  fabric_llpp1_arid_s_o(8)
       , fabric_llpp1_arid_s_o10                     =>  fabric_llpp1_arid_s_o(9)
       , fabric_llpp1_arid_s_o11                     =>  fabric_llpp1_arid_s_o(10)
       , fabric_llpp1_arid_s_o12                     =>  fabric_llpp1_arid_s_o(11)
       , fabric_llpp1_arlen_s_o1                     =>  fabric_llpp1_arlen_s_o(0)
       , fabric_llpp1_arlen_s_o2                     =>  fabric_llpp1_arlen_s_o(1)
       , fabric_llpp1_arlen_s_o3                     =>  fabric_llpp1_arlen_s_o(2)
       , fabric_llpp1_arlen_s_o4                     =>  fabric_llpp1_arlen_s_o(3)
       , fabric_llpp1_arlen_s_o5                     =>  fabric_llpp1_arlen_s_o(4)
       , fabric_llpp1_arlen_s_o6                     =>  fabric_llpp1_arlen_s_o(5)
       , fabric_llpp1_arlen_s_o7                     =>  fabric_llpp1_arlen_s_o(6)
       , fabric_llpp1_arlen_s_o8                     =>  fabric_llpp1_arlen_s_o(7)
       , fabric_llpp1_arlock_s_o                     =>  fabric_llpp1_arlock_s_o
       , fabric_llpp1_arprot_s_o1                    =>  fabric_llpp1_arprot_s_o(0)
       , fabric_llpp1_arprot_s_o2                    =>  fabric_llpp1_arprot_s_o(1)
       , fabric_llpp1_arprot_s_o3                    =>  fabric_llpp1_arprot_s_o(2)
       , fabric_llpp1_arqos_s1_o1                    =>  fabric_llpp1_arqos_s1_o(0)
       , fabric_llpp1_arqos_s1_o2                    =>  fabric_llpp1_arqos_s1_o(1)
       , fabric_llpp1_arqos_s1_o3                    =>  fabric_llpp1_arqos_s1_o(2)
       , fabric_llpp1_arqos_s1_o4                    =>  fabric_llpp1_arqos_s1_o(3)
       , fabric_llpp1_arsize_s_o1                    =>  fabric_llpp1_arsize_s_o(0)
       , fabric_llpp1_arsize_s_o2                    =>  fabric_llpp1_arsize_s_o(1)
       , fabric_llpp1_arsize_s_o3                    =>  fabric_llpp1_arsize_s_o(2)
       , fabric_llpp1_arvalid_s_o                    =>  fabric_llpp1_arvalid_s_o
       , fabric_llpp1_awaddr_s_o1                    =>  fabric_llpp1_awaddr_s_o(0)
       , fabric_llpp1_awaddr_s_o2                    =>  fabric_llpp1_awaddr_s_o(1)
       , fabric_llpp1_awaddr_s_o3                    =>  fabric_llpp1_awaddr_s_o(2)
       , fabric_llpp1_awaddr_s_o4                    =>  fabric_llpp1_awaddr_s_o(3)
       , fabric_llpp1_awaddr_s_o5                    =>  fabric_llpp1_awaddr_s_o(4)
       , fabric_llpp1_awaddr_s_o6                    =>  fabric_llpp1_awaddr_s_o(5)
       , fabric_llpp1_awaddr_s_o7                    =>  fabric_llpp1_awaddr_s_o(6)
       , fabric_llpp1_awaddr_s_o8                    =>  fabric_llpp1_awaddr_s_o(7)
       , fabric_llpp1_awaddr_s_o9                    =>  fabric_llpp1_awaddr_s_o(8)
       , fabric_llpp1_awaddr_s_o10                   =>  fabric_llpp1_awaddr_s_o(9)
       , fabric_llpp1_awaddr_s_o11                   =>  fabric_llpp1_awaddr_s_o(10)
       , fabric_llpp1_awaddr_s_o12                   =>  fabric_llpp1_awaddr_s_o(11)
       , fabric_llpp1_awaddr_s_o13                   =>  fabric_llpp1_awaddr_s_o(12)
       , fabric_llpp1_awaddr_s_o14                   =>  fabric_llpp1_awaddr_s_o(13)
       , fabric_llpp1_awaddr_s_o15                   =>  fabric_llpp1_awaddr_s_o(14)
       , fabric_llpp1_awaddr_s_o16                   =>  fabric_llpp1_awaddr_s_o(15)
       , fabric_llpp1_awaddr_s_o17                   =>  fabric_llpp1_awaddr_s_o(16)
       , fabric_llpp1_awaddr_s_o18                   =>  fabric_llpp1_awaddr_s_o(17)
       , fabric_llpp1_awaddr_s_o19                   =>  fabric_llpp1_awaddr_s_o(18)
       , fabric_llpp1_awaddr_s_o20                   =>  fabric_llpp1_awaddr_s_o(19)
       , fabric_llpp1_awaddr_s_o21                   =>  fabric_llpp1_awaddr_s_o(20)
       , fabric_llpp1_awaddr_s_o22                   =>  fabric_llpp1_awaddr_s_o(21)
       , fabric_llpp1_awaddr_s_o23                   =>  fabric_llpp1_awaddr_s_o(22)
       , fabric_llpp1_awaddr_s_o24                   =>  fabric_llpp1_awaddr_s_o(23)
       , fabric_llpp1_awaddr_s_o25                   =>  fabric_llpp1_awaddr_s_o(24)
       , fabric_llpp1_awaddr_s_o26                   =>  fabric_llpp1_awaddr_s_o(25)
       , fabric_llpp1_awaddr_s_o27                   =>  fabric_llpp1_awaddr_s_o(26)
       , fabric_llpp1_awaddr_s_o28                   =>  fabric_llpp1_awaddr_s_o(27)
       , fabric_llpp1_awaddr_s_o29                   =>  fabric_llpp1_awaddr_s_o(28)
       , fabric_llpp1_awaddr_s_o30                   =>  fabric_llpp1_awaddr_s_o(29)
       , fabric_llpp1_awaddr_s_o31                   =>  fabric_llpp1_awaddr_s_o(30)
       , fabric_llpp1_awaddr_s_o32                   =>  fabric_llpp1_awaddr_s_o(31)
       , fabric_llpp1_awburst_s_o1                   =>  fabric_llpp1_awburst_s_o(0)
       , fabric_llpp1_awburst_s_o2                   =>  fabric_llpp1_awburst_s_o(1)
       , fabric_llpp1_awcache_s_o1                   =>  fabric_llpp1_awcache_s_o(0)
       , fabric_llpp1_awcache_s_o2                   =>  fabric_llpp1_awcache_s_o(1)
       , fabric_llpp1_awcache_s_o3                   =>  fabric_llpp1_awcache_s_o(2)
       , fabric_llpp1_awcache_s_o4                   =>  fabric_llpp1_awcache_s_o(3)
       , fabric_llpp1_awid_s_o1                      =>  fabric_llpp1_awid_s_o(0)
       , fabric_llpp1_awid_s_o2                      =>  fabric_llpp1_awid_s_o(1)
       , fabric_llpp1_awid_s_o3                      =>  fabric_llpp1_awid_s_o(2)
       , fabric_llpp1_awid_s_o4                      =>  fabric_llpp1_awid_s_o(3)
       , fabric_llpp1_awid_s_o5                      =>  fabric_llpp1_awid_s_o(4)
       , fabric_llpp1_awid_s_o6                      =>  fabric_llpp1_awid_s_o(5)
       , fabric_llpp1_awid_s_o7                      =>  fabric_llpp1_awid_s_o(6)
       , fabric_llpp1_awid_s_o8                      =>  fabric_llpp1_awid_s_o(7)
       , fabric_llpp1_awid_s_o9                      =>  fabric_llpp1_awid_s_o(8)
       , fabric_llpp1_awid_s_o10                     =>  fabric_llpp1_awid_s_o(9)
       , fabric_llpp1_awid_s_o11                     =>  fabric_llpp1_awid_s_o(10)
       , fabric_llpp1_awid_s_o12                     =>  fabric_llpp1_awid_s_o(11)
       , fabric_llpp1_awlen_s_o1                     =>  fabric_llpp1_awlen_s_o(0)
       , fabric_llpp1_awlen_s_o2                     =>  fabric_llpp1_awlen_s_o(1)
       , fabric_llpp1_awlen_s_o3                     =>  fabric_llpp1_awlen_s_o(2)
       , fabric_llpp1_awlen_s_o4                     =>  fabric_llpp1_awlen_s_o(3)
       , fabric_llpp1_awlen_s_o5                     =>  fabric_llpp1_awlen_s_o(4)
       , fabric_llpp1_awlen_s_o6                     =>  fabric_llpp1_awlen_s_o(5)
       , fabric_llpp1_awlen_s_o7                     =>  fabric_llpp1_awlen_s_o(6)
       , fabric_llpp1_awlen_s_o8                     =>  fabric_llpp1_awlen_s_o(7)
       , fabric_llpp1_awlock_s_o                     =>  fabric_llpp1_awlock_s_o
       , fabric_llpp1_awprot_s_o1                    =>  fabric_llpp1_awprot_s_o(0)
       , fabric_llpp1_awprot_s_o2                    =>  fabric_llpp1_awprot_s_o(1)
       , fabric_llpp1_awprot_s_o3                    =>  fabric_llpp1_awprot_s_o(2)
       , fabric_llpp1_awqos_s_o1                     =>  fabric_llpp1_awqos_s_o(0)
       , fabric_llpp1_awqos_s_o2                     =>  fabric_llpp1_awqos_s_o(1)
       , fabric_llpp1_awqos_s_o3                     =>  fabric_llpp1_awqos_s_o(2)
       , fabric_llpp1_awqos_s_o4                     =>  fabric_llpp1_awqos_s_o(3)
       , fabric_llpp1_awsize_s_o1                    =>  fabric_llpp1_awsize_s_o(0)
       , fabric_llpp1_awsize_s_o2                    =>  fabric_llpp1_awsize_s_o(1)
       , fabric_llpp1_awsize_s_o3                    =>  fabric_llpp1_awsize_s_o(2)
       , fabric_llpp1_awvalid_s_o                    =>  fabric_llpp1_awvalid_s_o
       , fabric_llpp1_bready_s_o                     =>  fabric_llpp1_bready_s_o
       , fabric_llpp1_rready_s_o                     =>  fabric_llpp1_rready_s_o
       , fabric_llpp1_wdata_s_o1                     =>  fabric_llpp1_wdata_s_o(0)
       , fabric_llpp1_wdata_s_o2                     =>  fabric_llpp1_wdata_s_o(1)
       , fabric_llpp1_wdata_s_o3                     =>  fabric_llpp1_wdata_s_o(2)
       , fabric_llpp1_wdata_s_o4                     =>  fabric_llpp1_wdata_s_o(3)
       , fabric_llpp1_wdata_s_o5                     =>  fabric_llpp1_wdata_s_o(4)
       , fabric_llpp1_wdata_s_o6                     =>  fabric_llpp1_wdata_s_o(5)
       , fabric_llpp1_wdata_s_o7                     =>  fabric_llpp1_wdata_s_o(6)
       , fabric_llpp1_wdata_s_o8                     =>  fabric_llpp1_wdata_s_o(7)
       , fabric_llpp1_wdata_s_o9                     =>  fabric_llpp1_wdata_s_o(8)
       , fabric_llpp1_wdata_s_o10                    =>  fabric_llpp1_wdata_s_o(9)
       , fabric_llpp1_wdata_s_o11                    =>  fabric_llpp1_wdata_s_o(10)
       , fabric_llpp1_wdata_s_o12                    =>  fabric_llpp1_wdata_s_o(11)
       , fabric_llpp1_wdata_s_o13                    =>  fabric_llpp1_wdata_s_o(12)
       , fabric_llpp1_wdata_s_o14                    =>  fabric_llpp1_wdata_s_o(13)
       , fabric_llpp1_wdata_s_o15                    =>  fabric_llpp1_wdata_s_o(14)
       , fabric_llpp1_wdata_s_o16                    =>  fabric_llpp1_wdata_s_o(15)
       , fabric_llpp1_wdata_s_o17                    =>  fabric_llpp1_wdata_s_o(16)
       , fabric_llpp1_wdata_s_o18                    =>  fabric_llpp1_wdata_s_o(17)
       , fabric_llpp1_wdata_s_o19                    =>  fabric_llpp1_wdata_s_o(18)
       , fabric_llpp1_wdata_s_o20                    =>  fabric_llpp1_wdata_s_o(19)
       , fabric_llpp1_wdata_s_o21                    =>  fabric_llpp1_wdata_s_o(20)
       , fabric_llpp1_wdata_s_o22                    =>  fabric_llpp1_wdata_s_o(21)
       , fabric_llpp1_wdata_s_o23                    =>  fabric_llpp1_wdata_s_o(22)
       , fabric_llpp1_wdata_s_o24                    =>  fabric_llpp1_wdata_s_o(23)
       , fabric_llpp1_wdata_s_o25                    =>  fabric_llpp1_wdata_s_o(24)
       , fabric_llpp1_wdata_s_o26                    =>  fabric_llpp1_wdata_s_o(25)
       , fabric_llpp1_wdata_s_o27                    =>  fabric_llpp1_wdata_s_o(26)
       , fabric_llpp1_wdata_s_o28                    =>  fabric_llpp1_wdata_s_o(27)
       , fabric_llpp1_wdata_s_o29                    =>  fabric_llpp1_wdata_s_o(28)
       , fabric_llpp1_wdata_s_o30                    =>  fabric_llpp1_wdata_s_o(29)
       , fabric_llpp1_wdata_s_o31                    =>  fabric_llpp1_wdata_s_o(30)
       , fabric_llpp1_wdata_s_o32                    =>  fabric_llpp1_wdata_s_o(31)
       , fabric_llpp1_wlast_s_o                      =>  fabric_llpp1_wlast_s_o
       , fabric_llpp1_wstrb_s_o1                     =>  fabric_llpp1_wstrb_s_o(0)
       , fabric_llpp1_wstrb_s_o2                     =>  fabric_llpp1_wstrb_s_o(1)
       , fabric_llpp1_wstrb_s_o3                     =>  fabric_llpp1_wstrb_s_o(2)
       , fabric_llpp1_wstrb_s_o4                     =>  fabric_llpp1_wstrb_s_o(3)
       , fabric_llpp1_wvalid_s_o                     =>  fabric_llpp1_wvalid_s_o
       , fabric_llpp1_arready_s_i                    =>  fabric_llpp1_arready_s_i
       , fabric_llpp1_awready_s_i                    =>  fabric_llpp1_awready_s_i
       , fabric_llpp1_bid_s_i1                       =>  fabric_llpp1_bid_s_i(0)
       , fabric_llpp1_bid_s_i2                       =>  fabric_llpp1_bid_s_i(1)
       , fabric_llpp1_bid_s_i3                       =>  fabric_llpp1_bid_s_i(2)
       , fabric_llpp1_bid_s_i4                       =>  fabric_llpp1_bid_s_i(3)
       , fabric_llpp1_bid_s_i5                       =>  fabric_llpp1_bid_s_i(4)
       , fabric_llpp1_bid_s_i6                       =>  fabric_llpp1_bid_s_i(5)
       , fabric_llpp1_bid_s_i7                       =>  fabric_llpp1_bid_s_i(6)
       , fabric_llpp1_bid_s_i8                       =>  fabric_llpp1_bid_s_i(7)
       , fabric_llpp1_bid_s_i9                       =>  fabric_llpp1_bid_s_i(8)
       , fabric_llpp1_bid_s_i10                      =>  fabric_llpp1_bid_s_i(9)
       , fabric_llpp1_bid_s_i11                      =>  fabric_llpp1_bid_s_i(10)
       , fabric_llpp1_bid_s_i12                      =>  fabric_llpp1_bid_s_i(11)
       , fabric_llpp1_bresp_s_i1                     =>  fabric_llpp1_bresp_s_i(0)
       , fabric_llpp1_bresp_s_i2                     =>  fabric_llpp1_bresp_s_i(1)
       , fabric_llpp1_bvalid_s_i                     =>  fabric_llpp1_bvalid_s_i
       , fabric_llpp1_rdata_s_i1                     =>  fabric_llpp1_rdata_s_i(0)
       , fabric_llpp1_rdata_s_i2                     =>  fabric_llpp1_rdata_s_i(1)
       , fabric_llpp1_rdata_s_i3                     =>  fabric_llpp1_rdata_s_i(2)
       , fabric_llpp1_rdata_s_i4                     =>  fabric_llpp1_rdata_s_i(3)
       , fabric_llpp1_rdata_s_i5                     =>  fabric_llpp1_rdata_s_i(4)
       , fabric_llpp1_rdata_s_i6                     =>  fabric_llpp1_rdata_s_i(5)
       , fabric_llpp1_rdata_s_i7                     =>  fabric_llpp1_rdata_s_i(6)
       , fabric_llpp1_rdata_s_i8                     =>  fabric_llpp1_rdata_s_i(7)
       , fabric_llpp1_rdata_s_i9                     =>  fabric_llpp1_rdata_s_i(8)
       , fabric_llpp1_rdata_s_i10                    =>  fabric_llpp1_rdata_s_i(9)
       , fabric_llpp1_rdata_s_i11                    =>  fabric_llpp1_rdata_s_i(10)
       , fabric_llpp1_rdata_s_i12                    =>  fabric_llpp1_rdata_s_i(11)
       , fabric_llpp1_rdata_s_i13                    =>  fabric_llpp1_rdata_s_i(12)
       , fabric_llpp1_rdata_s_i14                    =>  fabric_llpp1_rdata_s_i(13)
       , fabric_llpp1_rdata_s_i15                    =>  fabric_llpp1_rdata_s_i(14)
       , fabric_llpp1_rdata_s_i16                    =>  fabric_llpp1_rdata_s_i(15)
       , fabric_llpp1_rdata_s_i17                    =>  fabric_llpp1_rdata_s_i(16)
       , fabric_llpp1_rdata_s_i18                    =>  fabric_llpp1_rdata_s_i(17)
       , fabric_llpp1_rdata_s_i19                    =>  fabric_llpp1_rdata_s_i(18)
       , fabric_llpp1_rdata_s_i20                    =>  fabric_llpp1_rdata_s_i(19)
       , fabric_llpp1_rdata_s_i21                    =>  fabric_llpp1_rdata_s_i(20)
       , fabric_llpp1_rdata_s_i22                    =>  fabric_llpp1_rdata_s_i(21)
       , fabric_llpp1_rdata_s_i23                    =>  fabric_llpp1_rdata_s_i(22)
       , fabric_llpp1_rdata_s_i24                    =>  fabric_llpp1_rdata_s_i(23)
       , fabric_llpp1_rdata_s_i25                    =>  fabric_llpp1_rdata_s_i(24)
       , fabric_llpp1_rdata_s_i26                    =>  fabric_llpp1_rdata_s_i(25)
       , fabric_llpp1_rdata_s_i27                    =>  fabric_llpp1_rdata_s_i(26)
       , fabric_llpp1_rdata_s_i28                    =>  fabric_llpp1_rdata_s_i(27)
       , fabric_llpp1_rdata_s_i29                    =>  fabric_llpp1_rdata_s_i(28)
       , fabric_llpp1_rdata_s_i30                    =>  fabric_llpp1_rdata_s_i(29)
       , fabric_llpp1_rdata_s_i31                    =>  fabric_llpp1_rdata_s_i(30)
       , fabric_llpp1_rdata_s_i32                    =>  fabric_llpp1_rdata_s_i(31)
       , fabric_llpp1_rid_s_i1                       =>  fabric_llpp1_rid_s_i(0)
       , fabric_llpp1_rid_s_i2                       =>  fabric_llpp1_rid_s_i(1)
       , fabric_llpp1_rid_s_i3                       =>  fabric_llpp1_rid_s_i(2)
       , fabric_llpp1_rid_s_i4                       =>  fabric_llpp1_rid_s_i(3)
       , fabric_llpp1_rid_s_i5                       =>  fabric_llpp1_rid_s_i(4)
       , fabric_llpp1_rid_s_i6                       =>  fabric_llpp1_rid_s_i(5)
       , fabric_llpp1_rid_s_i7                       =>  fabric_llpp1_rid_s_i(6)
       , fabric_llpp1_rid_s_i8                       =>  fabric_llpp1_rid_s_i(7)
       , fabric_llpp1_rid_s_i9                       =>  fabric_llpp1_rid_s_i(8)
       , fabric_llpp1_rid_s_i10                      =>  fabric_llpp1_rid_s_i(9)
       , fabric_llpp1_rid_s_i11                      =>  fabric_llpp1_rid_s_i(10)
       , fabric_llpp1_rid_s_i12                      =>  fabric_llpp1_rid_s_i(11)
       , fabric_llpp1_rlast_s_i                      =>  fabric_llpp1_rlast_s_i
       , fabric_llpp1_rresp_s_i1                     =>  fabric_llpp1_rresp_s_i(0)
       , fabric_llpp1_rresp_s_i2                     =>  fabric_llpp1_rresp_s_i(1)
       , fabric_llpp1_rvalid_s_i                     =>  fabric_llpp1_rvalid_s_i
       , fabric_llpp1_wready_s_i                     =>  fabric_llpp1_wready_s_i
       , fabric_llpp2_araddr_s_o1                    =>  fabric_llpp2_araddr_s_o(0)
       , fabric_llpp2_araddr_s_o2                    =>  fabric_llpp2_araddr_s_o(1)
       , fabric_llpp2_araddr_s_o3                    =>  fabric_llpp2_araddr_s_o(2)
       , fabric_llpp2_araddr_s_o4                    =>  fabric_llpp2_araddr_s_o(3)
       , fabric_llpp2_araddr_s_o5                    =>  fabric_llpp2_araddr_s_o(4)
       , fabric_llpp2_araddr_s_o6                    =>  fabric_llpp2_araddr_s_o(5)
       , fabric_llpp2_araddr_s_o7                    =>  fabric_llpp2_araddr_s_o(6)
       , fabric_llpp2_araddr_s_o8                    =>  fabric_llpp2_araddr_s_o(7)
       , fabric_llpp2_araddr_s_o9                    =>  fabric_llpp2_araddr_s_o(8)
       , fabric_llpp2_araddr_s_o10                   =>  fabric_llpp2_araddr_s_o(9)
       , fabric_llpp2_araddr_s_o11                   =>  fabric_llpp2_araddr_s_o(10)
       , fabric_llpp2_araddr_s_o12                   =>  fabric_llpp2_araddr_s_o(11)
       , fabric_llpp2_araddr_s_o13                   =>  fabric_llpp2_araddr_s_o(12)
       , fabric_llpp2_araddr_s_o14                   =>  fabric_llpp2_araddr_s_o(13)
       , fabric_llpp2_araddr_s_o15                   =>  fabric_llpp2_araddr_s_o(14)
       , fabric_llpp2_araddr_s_o16                   =>  fabric_llpp2_araddr_s_o(15)
       , fabric_llpp2_araddr_s_o17                   =>  fabric_llpp2_araddr_s_o(16)
       , fabric_llpp2_araddr_s_o18                   =>  fabric_llpp2_araddr_s_o(17)
       , fabric_llpp2_araddr_s_o19                   =>  fabric_llpp2_araddr_s_o(18)
       , fabric_llpp2_araddr_s_o20                   =>  fabric_llpp2_araddr_s_o(19)
       , fabric_llpp2_araddr_s_o21                   =>  fabric_llpp2_araddr_s_o(20)
       , fabric_llpp2_araddr_s_o22                   =>  fabric_llpp2_araddr_s_o(21)
       , fabric_llpp2_araddr_s_o23                   =>  fabric_llpp2_araddr_s_o(22)
       , fabric_llpp2_araddr_s_o24                   =>  fabric_llpp2_araddr_s_o(23)
       , fabric_llpp2_araddr_s_o25                   =>  fabric_llpp2_araddr_s_o(24)
       , fabric_llpp2_araddr_s_o26                   =>  fabric_llpp2_araddr_s_o(25)
       , fabric_llpp2_araddr_s_o27                   =>  fabric_llpp2_araddr_s_o(26)
       , fabric_llpp2_araddr_s_o28                   =>  fabric_llpp2_araddr_s_o(27)
       , fabric_llpp2_araddr_s_o29                   =>  fabric_llpp2_araddr_s_o(28)
       , fabric_llpp2_araddr_s_o30                   =>  fabric_llpp2_araddr_s_o(29)
       , fabric_llpp2_araddr_s_o31                   =>  fabric_llpp2_araddr_s_o(30)
       , fabric_llpp2_araddr_s_o32                   =>  fabric_llpp2_araddr_s_o(31)
       , fabric_llpp2_arburst_s_o1                   =>  fabric_llpp2_arburst_s_o(0)
       , fabric_llpp2_arburst_s_o2                   =>  fabric_llpp2_arburst_s_o(1)
       , fabric_llpp2_arcache_s_o1                   =>  fabric_llpp2_arcache_s_o(0)
       , fabric_llpp2_arcache_s_o2                   =>  fabric_llpp2_arcache_s_o(1)
       , fabric_llpp2_arcache_s_o3                   =>  fabric_llpp2_arcache_s_o(2)
       , fabric_llpp2_arcache_s_o4                   =>  fabric_llpp2_arcache_s_o(3)
       , fabric_llpp2_arid_s_o1                      =>  fabric_llpp2_arid_s_o(0)
       , fabric_llpp2_arid_s_o2                      =>  fabric_llpp2_arid_s_o(1)
       , fabric_llpp2_arid_s_o3                      =>  fabric_llpp2_arid_s_o(2)
       , fabric_llpp2_arid_s_o4                      =>  fabric_llpp2_arid_s_o(3)
       , fabric_llpp2_arid_s_o5                      =>  fabric_llpp2_arid_s_o(4)
       , fabric_llpp2_arid_s_o6                      =>  fabric_llpp2_arid_s_o(5)
       , fabric_llpp2_arid_s_o7                      =>  fabric_llpp2_arid_s_o(6)
       , fabric_llpp2_arid_s_o8                      =>  fabric_llpp2_arid_s_o(7)
       , fabric_llpp2_arid_s_o9                      =>  fabric_llpp2_arid_s_o(8)
       , fabric_llpp2_arid_s_o10                     =>  fabric_llpp2_arid_s_o(9)
       , fabric_llpp2_arid_s_o11                     =>  fabric_llpp2_arid_s_o(10)
       , fabric_llpp2_arid_s_o12                     =>  fabric_llpp2_arid_s_o(11)
       , fabric_llpp2_arlen_s_o1                     =>  fabric_llpp2_arlen_s_o(0)
       , fabric_llpp2_arlen_s_o2                     =>  fabric_llpp2_arlen_s_o(1)
       , fabric_llpp2_arlen_s_o3                     =>  fabric_llpp2_arlen_s_o(2)
       , fabric_llpp2_arlen_s_o4                     =>  fabric_llpp2_arlen_s_o(3)
       , fabric_llpp2_arlen_s_o5                     =>  fabric_llpp2_arlen_s_o(4)
       , fabric_llpp2_arlen_s_o6                     =>  fabric_llpp2_arlen_s_o(5)
       , fabric_llpp2_arlen_s_o7                     =>  fabric_llpp2_arlen_s_o(6)
       , fabric_llpp2_arlen_s_o8                     =>  fabric_llpp2_arlen_s_o(7)
       , fabric_llpp2_arlock_s_o                     =>  fabric_llpp2_arlock_s_o
       , fabric_llpp2_arprot_s_o1                    =>  fabric_llpp2_arprot_s_o(0)
       , fabric_llpp2_arprot_s_o2                    =>  fabric_llpp2_arprot_s_o(1)
       , fabric_llpp2_arprot_s_o3                    =>  fabric_llpp2_arprot_s_o(2)
       , fabric_llpp2_arqos_s_o1                     =>  fabric_llpp2_arqos_s_o(0)
       , fabric_llpp2_arqos_s_o2                     =>  fabric_llpp2_arqos_s_o(1)
       , fabric_llpp2_arqos_s_o3                     =>  fabric_llpp2_arqos_s_o(2)
       , fabric_llpp2_arqos_s_o4                     =>  fabric_llpp2_arqos_s_o(3)
       , fabric_llpp2_arsize_s_o1                    =>  fabric_llpp2_arsize_s_o(0)
       , fabric_llpp2_arsize_s_o2                    =>  fabric_llpp2_arsize_s_o(1)
       , fabric_llpp2_arsize_s_o3                    =>  fabric_llpp2_arsize_s_o(2)
       , fabric_llpp2_arvalid_s_o                    =>  fabric_llpp2_arvalid_s_o
       , fabric_llpp2_awaddr_s_o1                    =>  fabric_llpp2_awaddr_s_o(0)
       , fabric_llpp2_awaddr_s_o2                    =>  fabric_llpp2_awaddr_s_o(1)
       , fabric_llpp2_awaddr_s_o3                    =>  fabric_llpp2_awaddr_s_o(2)
       , fabric_llpp2_awaddr_s_o4                    =>  fabric_llpp2_awaddr_s_o(3)
       , fabric_llpp2_awaddr_s_o5                    =>  fabric_llpp2_awaddr_s_o(4)
       , fabric_llpp2_awaddr_s_o6                    =>  fabric_llpp2_awaddr_s_o(5)
       , fabric_llpp2_awaddr_s_o7                    =>  fabric_llpp2_awaddr_s_o(6)
       , fabric_llpp2_awaddr_s_o8                    =>  fabric_llpp2_awaddr_s_o(7)
       , fabric_llpp2_awaddr_s_o9                    =>  fabric_llpp2_awaddr_s_o(8)
       , fabric_llpp2_awaddr_s_o10                   =>  fabric_llpp2_awaddr_s_o(9)
       , fabric_llpp2_awaddr_s_o11                   =>  fabric_llpp2_awaddr_s_o(10)
       , fabric_llpp2_awaddr_s_o12                   =>  fabric_llpp2_awaddr_s_o(11)
       , fabric_llpp2_awaddr_s_o13                   =>  fabric_llpp2_awaddr_s_o(12)
       , fabric_llpp2_awaddr_s_o14                   =>  fabric_llpp2_awaddr_s_o(13)
       , fabric_llpp2_awaddr_s_o15                   =>  fabric_llpp2_awaddr_s_o(14)
       , fabric_llpp2_awaddr_s_o16                   =>  fabric_llpp2_awaddr_s_o(15)
       , fabric_llpp2_awaddr_s_o17                   =>  fabric_llpp2_awaddr_s_o(16)
       , fabric_llpp2_awaddr_s_o18                   =>  fabric_llpp2_awaddr_s_o(17)
       , fabric_llpp2_awaddr_s_o19                   =>  fabric_llpp2_awaddr_s_o(18)
       , fabric_llpp2_awaddr_s_o20                   =>  fabric_llpp2_awaddr_s_o(19)
       , fabric_llpp2_awaddr_s_o21                   =>  fabric_llpp2_awaddr_s_o(20)
       , fabric_llpp2_awaddr_s_o22                   =>  fabric_llpp2_awaddr_s_o(21)
       , fabric_llpp2_awaddr_s_o23                   =>  fabric_llpp2_awaddr_s_o(22)
       , fabric_llpp2_awaddr_s_o24                   =>  fabric_llpp2_awaddr_s_o(23)
       , fabric_llpp2_awaddr_s_o25                   =>  fabric_llpp2_awaddr_s_o(24)
       , fabric_llpp2_awaddr_s_o26                   =>  fabric_llpp2_awaddr_s_o(25)
       , fabric_llpp2_awaddr_s_o27                   =>  fabric_llpp2_awaddr_s_o(26)
       , fabric_llpp2_awaddr_s_o28                   =>  fabric_llpp2_awaddr_s_o(27)
       , fabric_llpp2_awaddr_s_o29                   =>  fabric_llpp2_awaddr_s_o(28)
       , fabric_llpp2_awaddr_s_o30                   =>  fabric_llpp2_awaddr_s_o(29)
       , fabric_llpp2_awaddr_s_o31                   =>  fabric_llpp2_awaddr_s_o(30)
       , fabric_llpp2_awaddr_s_o32                   =>  fabric_llpp2_awaddr_s_o(31)
       , fabric_llpp2_awburst_s_o1                   =>  fabric_llpp2_awburst_s_o(0)
       , fabric_llpp2_awburst_s_o2                   =>  fabric_llpp2_awburst_s_o(1)
       , fabric_llpp2_awcache_s_o1                   =>  fabric_llpp2_awcache_s_o(0)
       , fabric_llpp2_awcache_s_o2                   =>  fabric_llpp2_awcache_s_o(1)
       , fabric_llpp2_awcache_s_o3                   =>  fabric_llpp2_awcache_s_o(2)
       , fabric_llpp2_awcache_s_o4                   =>  fabric_llpp2_awcache_s_o(3)
       , fabric_llpp2_awid_s_o1                      =>  fabric_llpp2_awid_s_o(0)
       , fabric_llpp2_awid_s_o2                      =>  fabric_llpp2_awid_s_o(1)
       , fabric_llpp2_awid_s_o3                      =>  fabric_llpp2_awid_s_o(2)
       , fabric_llpp2_awid_s_o4                      =>  fabric_llpp2_awid_s_o(3)
       , fabric_llpp2_awid_s_o5                      =>  fabric_llpp2_awid_s_o(4)
       , fabric_llpp2_awid_s_o6                      =>  fabric_llpp2_awid_s_o(5)
       , fabric_llpp2_awid_s_o7                      =>  fabric_llpp2_awid_s_o(6)
       , fabric_llpp2_awid_s_o8                      =>  fabric_llpp2_awid_s_o(7)
       , fabric_llpp2_awid_s_o9                      =>  fabric_llpp2_awid_s_o(8)
       , fabric_llpp2_awid_s_o10                     =>  fabric_llpp2_awid_s_o(9)
       , fabric_llpp2_awid_s_o11                     =>  fabric_llpp2_awid_s_o(10)
       , fabric_llpp2_awid_s_o12                     =>  fabric_llpp2_awid_s_o(11)
       , fabric_llpp2_awlen_s_o1                     =>  fabric_llpp2_awlen_s_o(0)
       , fabric_llpp2_awlen_s_o2                     =>  fabric_llpp2_awlen_s_o(1)
       , fabric_llpp2_awlen_s_o3                     =>  fabric_llpp2_awlen_s_o(2)
       , fabric_llpp2_awlen_s_o4                     =>  fabric_llpp2_awlen_s_o(3)
       , fabric_llpp2_awlen_s_o5                     =>  fabric_llpp2_awlen_s_o(4)
       , fabric_llpp2_awlen_s_o6                     =>  fabric_llpp2_awlen_s_o(5)
       , fabric_llpp2_awlen_s_o7                     =>  fabric_llpp2_awlen_s_o(6)
       , fabric_llpp2_awlen_s_o8                     =>  fabric_llpp2_awlen_s_o(7)
       , fabric_llpp2_awlock_s_o                     =>  fabric_llpp2_awlock_s_o
       , fabric_llpp2_awprot_s_o1                    =>  fabric_llpp2_awprot_s_o(0)
       , fabric_llpp2_awprot_s_o2                    =>  fabric_llpp2_awprot_s_o(1)
       , fabric_llpp2_awprot_s_o3                    =>  fabric_llpp2_awprot_s_o(2)
       , fabric_llpp2_awqos_s_o1                     =>  fabric_llpp2_awqos_s_o(0)
       , fabric_llpp2_awqos_s_o2                     =>  fabric_llpp2_awqos_s_o(1)
       , fabric_llpp2_awqos_s_o3                     =>  fabric_llpp2_awqos_s_o(2)
       , fabric_llpp2_awqos_s_o4                     =>  fabric_llpp2_awqos_s_o(3)
       , fabric_llpp2_awsize_s_o1                    =>  fabric_llpp2_awsize_s_o(0)
       , fabric_llpp2_awsize_s_o2                    =>  fabric_llpp2_awsize_s_o(1)
       , fabric_llpp2_awsize_s_o3                    =>  fabric_llpp2_awsize_s_o(2)
       , fabric_llpp2_awvalid_s_o                    =>  fabric_llpp2_awvalid_s_o
       , fabric_llpp2_bready_s_o                     =>  fabric_llpp2_bready_s_o
       , fabric_llpp2_rready_s_o                     =>  fabric_llpp2_rready_s_o
       , fabric_llpp2_wdata_s_o1                     =>  fabric_llpp2_wdata_s_o(0)
       , fabric_llpp2_wdata_s_o2                     =>  fabric_llpp2_wdata_s_o(1)
       , fabric_llpp2_wdata_s_o3                     =>  fabric_llpp2_wdata_s_o(2)
       , fabric_llpp2_wdata_s_o4                     =>  fabric_llpp2_wdata_s_o(3)
       , fabric_llpp2_wdata_s_o5                     =>  fabric_llpp2_wdata_s_o(4)
       , fabric_llpp2_wdata_s_o6                     =>  fabric_llpp2_wdata_s_o(5)
       , fabric_llpp2_wdata_s_o7                     =>  fabric_llpp2_wdata_s_o(6)
       , fabric_llpp2_wdata_s_o8                     =>  fabric_llpp2_wdata_s_o(7)
       , fabric_llpp2_wdata_s_o9                     =>  fabric_llpp2_wdata_s_o(8)
       , fabric_llpp2_wdata_s_o10                    =>  fabric_llpp2_wdata_s_o(9)
       , fabric_llpp2_wdata_s_o11                    =>  fabric_llpp2_wdata_s_o(10)
       , fabric_llpp2_wdata_s_o12                    =>  fabric_llpp2_wdata_s_o(11)
       , fabric_llpp2_wdata_s_o13                    =>  fabric_llpp2_wdata_s_o(12)
       , fabric_llpp2_wdata_s_o14                    =>  fabric_llpp2_wdata_s_o(13)
       , fabric_llpp2_wdata_s_o15                    =>  fabric_llpp2_wdata_s_o(14)
       , fabric_llpp2_wdata_s_o16                    =>  fabric_llpp2_wdata_s_o(15)
       , fabric_llpp2_wdata_s_o17                    =>  fabric_llpp2_wdata_s_o(16)
       , fabric_llpp2_wdata_s_o18                    =>  fabric_llpp2_wdata_s_o(17)
       , fabric_llpp2_wdata_s_o19                    =>  fabric_llpp2_wdata_s_o(18)
       , fabric_llpp2_wdata_s_o20                    =>  fabric_llpp2_wdata_s_o(19)
       , fabric_llpp2_wdata_s_o21                    =>  fabric_llpp2_wdata_s_o(20)
       , fabric_llpp2_wdata_s_o22                    =>  fabric_llpp2_wdata_s_o(21)
       , fabric_llpp2_wdata_s_o23                    =>  fabric_llpp2_wdata_s_o(22)
       , fabric_llpp2_wdata_s_o24                    =>  fabric_llpp2_wdata_s_o(23)
       , fabric_llpp2_wdata_s_o25                    =>  fabric_llpp2_wdata_s_o(24)
       , fabric_llpp2_wdata_s_o26                    =>  fabric_llpp2_wdata_s_o(25)
       , fabric_llpp2_wdata_s_o27                    =>  fabric_llpp2_wdata_s_o(26)
       , fabric_llpp2_wdata_s_o28                    =>  fabric_llpp2_wdata_s_o(27)
       , fabric_llpp2_wdata_s_o29                    =>  fabric_llpp2_wdata_s_o(28)
       , fabric_llpp2_wdata_s_o30                    =>  fabric_llpp2_wdata_s_o(29)
       , fabric_llpp2_wdata_s_o31                    =>  fabric_llpp2_wdata_s_o(30)
       , fabric_llpp2_wdata_s_o32                    =>  fabric_llpp2_wdata_s_o(31)
       , fabric_llpp2_wlast_s_o                      =>  fabric_llpp2_wlast_s_o
       , fabric_llpp2_wstrb_s_o1                     =>  fabric_llpp2_wstrb_s_o(0)
       , fabric_llpp2_wstrb_s_o2                     =>  fabric_llpp2_wstrb_s_o(1)
       , fabric_llpp2_wstrb_s_o3                     =>  fabric_llpp2_wstrb_s_o(2)
       , fabric_llpp2_wstrb_s_o4                     =>  fabric_llpp2_wstrb_s_o(3)
       , fabric_llpp2_wvalid_s_o                     =>  fabric_llpp2_wvalid_s_o
       , fabric_llpp2_arready_s_i                    =>  fabric_llpp2_arready_s_i
       , fabric_llpp2_awready_s_i                    =>  fabric_llpp2_awready_s_i
       , fabric_llpp2_bid_s_i1                       =>  fabric_llpp2_bid_s_i(0)
       , fabric_llpp2_bid_s_i2                       =>  fabric_llpp2_bid_s_i(1)
       , fabric_llpp2_bid_s_i3                       =>  fabric_llpp2_bid_s_i(2)
       , fabric_llpp2_bid_s_i4                       =>  fabric_llpp2_bid_s_i(3)
       , fabric_llpp2_bid_s_i5                       =>  fabric_llpp2_bid_s_i(4)
       , fabric_llpp2_bid_s_i6                       =>  fabric_llpp2_bid_s_i(5)
       , fabric_llpp2_bid_s_i7                       =>  fabric_llpp2_bid_s_i(6)
       , fabric_llpp2_bid_s_i8                       =>  fabric_llpp2_bid_s_i(7)
       , fabric_llpp2_bid_s_i9                       =>  fabric_llpp2_bid_s_i(8)
       , fabric_llpp2_bid_s_i10                      =>  fabric_llpp2_bid_s_i(9)
       , fabric_llpp2_bid_s_i11                      =>  fabric_llpp2_bid_s_i(10)
       , fabric_llpp2_bid_s_i12                      =>  fabric_llpp2_bid_s_i(11)
       , fabric_llpp2_bresp_s_i1                     =>  fabric_llpp2_bresp_s_i(0)
       , fabric_llpp2_bresp_s_i2                     =>  fabric_llpp2_bresp_s_i(1)
       , fabric_llpp2_bvalid_s_i                     =>  fabric_llpp2_bvalid_s_i
       , fabric_llpp2_rdata_s_i1                     =>  fabric_llpp2_rdata_s_i(0)
       , fabric_llpp2_rdata_s_i2                     =>  fabric_llpp2_rdata_s_i(1)
       , fabric_llpp2_rdata_s_i3                     =>  fabric_llpp2_rdata_s_i(2)
       , fabric_llpp2_rdata_s_i4                     =>  fabric_llpp2_rdata_s_i(3)
       , fabric_llpp2_rdata_s_i5                     =>  fabric_llpp2_rdata_s_i(4)
       , fabric_llpp2_rdata_s_i6                     =>  fabric_llpp2_rdata_s_i(5)
       , fabric_llpp2_rdata_s_i7                     =>  fabric_llpp2_rdata_s_i(6)
       , fabric_llpp2_rdata_s_i8                     =>  fabric_llpp2_rdata_s_i(7)
       , fabric_llpp2_rdata_s_i9                     =>  fabric_llpp2_rdata_s_i(8)
       , fabric_llpp2_rdata_s_i10                    =>  fabric_llpp2_rdata_s_i(9)
       , fabric_llpp2_rdata_s_i11                    =>  fabric_llpp2_rdata_s_i(10)
       , fabric_llpp2_rdata_s_i12                    =>  fabric_llpp2_rdata_s_i(11)
       , fabric_llpp2_rdata_s_i13                    =>  fabric_llpp2_rdata_s_i(12)
       , fabric_llpp2_rdata_s_i14                    =>  fabric_llpp2_rdata_s_i(13)
       , fabric_llpp2_rdata_s_i15                    =>  fabric_llpp2_rdata_s_i(14)
       , fabric_llpp2_rdata_s_i16                    =>  fabric_llpp2_rdata_s_i(15)
       , fabric_llpp2_rdata_s_i17                    =>  fabric_llpp2_rdata_s_i(16)
       , fabric_llpp2_rdata_s_i18                    =>  fabric_llpp2_rdata_s_i(17)
       , fabric_llpp2_rdata_s_i19                    =>  fabric_llpp2_rdata_s_i(18)
       , fabric_llpp2_rdata_s_i20                    =>  fabric_llpp2_rdata_s_i(19)
       , fabric_llpp2_rdata_s_i21                    =>  fabric_llpp2_rdata_s_i(20)
       , fabric_llpp2_rdata_s_i22                    =>  fabric_llpp2_rdata_s_i(21)
       , fabric_llpp2_rdata_s_i23                    =>  fabric_llpp2_rdata_s_i(22)
       , fabric_llpp2_rdata_s_i24                    =>  fabric_llpp2_rdata_s_i(23)
       , fabric_llpp2_rdata_s_i25                    =>  fabric_llpp2_rdata_s_i(24)
       , fabric_llpp2_rdata_s_i26                    =>  fabric_llpp2_rdata_s_i(25)
       , fabric_llpp2_rdata_s_i27                    =>  fabric_llpp2_rdata_s_i(26)
       , fabric_llpp2_rdata_s_i28                    =>  fabric_llpp2_rdata_s_i(27)
       , fabric_llpp2_rdata_s_i29                    =>  fabric_llpp2_rdata_s_i(28)
       , fabric_llpp2_rdata_s_i30                    =>  fabric_llpp2_rdata_s_i(29)
       , fabric_llpp2_rdata_s_i31                    =>  fabric_llpp2_rdata_s_i(30)
       , fabric_llpp2_rdata_s_i32                    =>  fabric_llpp2_rdata_s_i(31)
       , fabric_llpp2_rid_s_i1                       =>  fabric_llpp2_rid_s_i(0)
       , fabric_llpp2_rid_s_i2                       =>  fabric_llpp2_rid_s_i(1)
       , fabric_llpp2_rid_s_i3                       =>  fabric_llpp2_rid_s_i(2)
       , fabric_llpp2_rid_s_i4                       =>  fabric_llpp2_rid_s_i(3)
       , fabric_llpp2_rid_s_i5                       =>  fabric_llpp2_rid_s_i(4)
       , fabric_llpp2_rid_s_i6                       =>  fabric_llpp2_rid_s_i(5)
       , fabric_llpp2_rid_s_i7                       =>  fabric_llpp2_rid_s_i(6)
       , fabric_llpp2_rid_s_i8                       =>  fabric_llpp2_rid_s_i(7)
       , fabric_llpp2_rid_s_i9                       =>  fabric_llpp2_rid_s_i(8)
       , fabric_llpp2_rid_s_i10                      =>  fabric_llpp2_rid_s_i(9)
       , fabric_llpp2_rid_s_i11                      =>  fabric_llpp2_rid_s_i(10)
       , fabric_llpp2_rid_s_i12                      =>  fabric_llpp2_rid_s_i(11)
       , fabric_llpp2_rlast_s_i                      =>  fabric_llpp2_rlast_s_i
       , fabric_llpp2_rresp_s_i1                     =>  fabric_llpp2_rresp_s_i(0)
       , fabric_llpp2_rresp_s_i2                     =>  fabric_llpp2_rresp_s_i(1)
       , fabric_llpp2_rvalid_s_i                     =>  fabric_llpp2_rvalid_s_i
       , fabric_llpp2_wready_s_i                     =>  fabric_llpp2_wready_s_i
       , fabric_llpp3_araddr_s_o1                    =>  fabric_llpp3_araddr_s_o(0)
       , fabric_llpp3_araddr_s_o2                    =>  fabric_llpp3_araddr_s_o(1)
       , fabric_llpp3_araddr_s_o3                    =>  fabric_llpp3_araddr_s_o(2)
       , fabric_llpp3_araddr_s_o4                    =>  fabric_llpp3_araddr_s_o(3)
       , fabric_llpp3_araddr_s_o5                    =>  fabric_llpp3_araddr_s_o(4)
       , fabric_llpp3_araddr_s_o6                    =>  fabric_llpp3_araddr_s_o(5)
       , fabric_llpp3_araddr_s_o7                    =>  fabric_llpp3_araddr_s_o(6)
       , fabric_llpp3_araddr_s_o8                    =>  fabric_llpp3_araddr_s_o(7)
       , fabric_llpp3_araddr_s_o9                    =>  fabric_llpp3_araddr_s_o(8)
       , fabric_llpp3_araddr_s_o10                   =>  fabric_llpp3_araddr_s_o(9)
       , fabric_llpp3_araddr_s_o11                   =>  fabric_llpp3_araddr_s_o(10)
       , fabric_llpp3_araddr_s_o12                   =>  fabric_llpp3_araddr_s_o(11)
       , fabric_llpp3_araddr_s_o13                   =>  fabric_llpp3_araddr_s_o(12)
       , fabric_llpp3_araddr_s_o14                   =>  fabric_llpp3_araddr_s_o(13)
       , fabric_llpp3_araddr_s_o15                   =>  fabric_llpp3_araddr_s_o(14)
       , fabric_llpp3_araddr_s_o16                   =>  fabric_llpp3_araddr_s_o(15)
       , fabric_llpp3_araddr_s_o17                   =>  fabric_llpp3_araddr_s_o(16)
       , fabric_llpp3_araddr_s_o18                   =>  fabric_llpp3_araddr_s_o(17)
       , fabric_llpp3_araddr_s_o19                   =>  fabric_llpp3_araddr_s_o(18)
       , fabric_llpp3_araddr_s_o20                   =>  fabric_llpp3_araddr_s_o(19)
       , fabric_llpp3_araddr_s_o21                   =>  fabric_llpp3_araddr_s_o(20)
       , fabric_llpp3_araddr_s_o22                   =>  fabric_llpp3_araddr_s_o(21)
       , fabric_llpp3_araddr_s_o23                   =>  fabric_llpp3_araddr_s_o(22)
       , fabric_llpp3_araddr_s_o24                   =>  fabric_llpp3_araddr_s_o(23)
       , fabric_llpp3_araddr_s_o25                   =>  fabric_llpp3_araddr_s_o(24)
       , fabric_llpp3_araddr_s_o26                   =>  fabric_llpp3_araddr_s_o(25)
       , fabric_llpp3_araddr_s_o27                   =>  fabric_llpp3_araddr_s_o(26)
       , fabric_llpp3_araddr_s_o28                   =>  fabric_llpp3_araddr_s_o(27)
       , fabric_llpp3_araddr_s_o29                   =>  fabric_llpp3_araddr_s_o(28)
       , fabric_llpp3_araddr_s_o30                   =>  fabric_llpp3_araddr_s_o(29)
       , fabric_llpp3_araddr_s_o31                   =>  fabric_llpp3_araddr_s_o(30)
       , fabric_llpp3_araddr_s_o32                   =>  fabric_llpp3_araddr_s_o(31)
       , fabric_llpp3_arburst_s_o1                   =>  fabric_llpp3_arburst_s_o(0)
       , fabric_llpp3_arburst_s_o2                   =>  fabric_llpp3_arburst_s_o(1)
       , fabric_llpp3_arcache_s_o1                   =>  fabric_llpp3_arcache_s_o(0)
       , fabric_llpp3_arcache_s_o2                   =>  fabric_llpp3_arcache_s_o(1)
       , fabric_llpp3_arcache_s_o3                   =>  fabric_llpp3_arcache_s_o(2)
       , fabric_llpp3_arcache_s_o4                   =>  fabric_llpp3_arcache_s_o(3)
       , fabric_llpp3_arid_s_o1                      =>  fabric_llpp3_arid_s_o(0)
       , fabric_llpp3_arid_s_o2                      =>  fabric_llpp3_arid_s_o(1)
       , fabric_llpp3_arid_s_o3                      =>  fabric_llpp3_arid_s_o(2)
       , fabric_llpp3_arid_s_o4                      =>  fabric_llpp3_arid_s_o(3)
       , fabric_llpp3_arid_s_o5                      =>  fabric_llpp3_arid_s_o(4)
       , fabric_llpp3_arid_s_o6                      =>  fabric_llpp3_arid_s_o(5)
       , fabric_llpp3_arid_s_o7                      =>  fabric_llpp3_arid_s_o(6)
       , fabric_llpp3_arid_s_o8                      =>  fabric_llpp3_arid_s_o(7)
       , fabric_llpp3_arid_s_o9                      =>  fabric_llpp3_arid_s_o(8)
       , fabric_llpp3_arid_s_o10                     =>  fabric_llpp3_arid_s_o(9)
       , fabric_llpp3_arid_s_o11                     =>  fabric_llpp3_arid_s_o(10)
       , fabric_llpp3_arid_s_o12                     =>  fabric_llpp3_arid_s_o(11)
       , fabric_llpp3_arlen_s_o1                     =>  fabric_llpp3_arlen_s_o(0)
       , fabric_llpp3_arlen_s_o2                     =>  fabric_llpp3_arlen_s_o(1)
       , fabric_llpp3_arlen_s_o3                     =>  fabric_llpp3_arlen_s_o(2)
       , fabric_llpp3_arlen_s_o4                     =>  fabric_llpp3_arlen_s_o(3)
       , fabric_llpp3_arlen_s_o5                     =>  fabric_llpp3_arlen_s_o(4)
       , fabric_llpp3_arlen_s_o6                     =>  fabric_llpp3_arlen_s_o(5)
       , fabric_llpp3_arlen_s_o7                     =>  fabric_llpp3_arlen_s_o(6)
       , fabric_llpp3_arlen_s_o8                     =>  fabric_llpp3_arlen_s_o(7)
       , fabric_llpp3_arlock_s_o                     =>  fabric_llpp3_arlock_s_o
       , fabric_llpp3_arprot_s_o1                    =>  fabric_llpp3_arprot_s_o(0)
       , fabric_llpp3_arprot_s_o2                    =>  fabric_llpp3_arprot_s_o(1)
       , fabric_llpp3_arprot_s_o3                    =>  fabric_llpp3_arprot_s_o(2)
       , fabric_llpp3_arqos_s_o1                     =>  fabric_llpp3_arqos_s_o(0)
       , fabric_llpp3_arqos_s_o2                     =>  fabric_llpp3_arqos_s_o(1)
       , fabric_llpp3_arqos_s_o3                     =>  fabric_llpp3_arqos_s_o(2)
       , fabric_llpp3_arqos_s_o4                     =>  fabric_llpp3_arqos_s_o(3)
       , fabric_llpp3_arsize_s_o1                    =>  fabric_llpp3_arsize_s_o(0)
       , fabric_llpp3_arsize_s_o2                    =>  fabric_llpp3_arsize_s_o(1)
       , fabric_llpp3_arsize_s_o3                    =>  fabric_llpp3_arsize_s_o(2)
       , fabric_llpp3_arvalid_s_o                    =>  fabric_llpp3_arvalid_s_o
       , fabric_llpp3_awaddr_s_o1                    =>  fabric_llpp3_awaddr_s_o(0)
       , fabric_llpp3_awaddr_s_o2                    =>  fabric_llpp3_awaddr_s_o(1)
       , fabric_llpp3_awaddr_s_o3                    =>  fabric_llpp3_awaddr_s_o(2)
       , fabric_llpp3_awaddr_s_o4                    =>  fabric_llpp3_awaddr_s_o(3)
       , fabric_llpp3_awaddr_s_o5                    =>  fabric_llpp3_awaddr_s_o(4)
       , fabric_llpp3_awaddr_s_o6                    =>  fabric_llpp3_awaddr_s_o(5)
       , fabric_llpp3_awaddr_s_o7                    =>  fabric_llpp3_awaddr_s_o(6)
       , fabric_llpp3_awaddr_s_o8                    =>  fabric_llpp3_awaddr_s_o(7)
       , fabric_llpp3_awaddr_s_o9                    =>  fabric_llpp3_awaddr_s_o(8)
       , fabric_llpp3_awaddr_s_o10                   =>  fabric_llpp3_awaddr_s_o(9)
       , fabric_llpp3_awaddr_s_o11                   =>  fabric_llpp3_awaddr_s_o(10)
       , fabric_llpp3_awaddr_s_o12                   =>  fabric_llpp3_awaddr_s_o(11)
       , fabric_llpp3_awaddr_s_o13                   =>  fabric_llpp3_awaddr_s_o(12)
       , fabric_llpp3_awaddr_s_o14                   =>  fabric_llpp3_awaddr_s_o(13)
       , fabric_llpp3_awaddr_s_o15                   =>  fabric_llpp3_awaddr_s_o(14)
       , fabric_llpp3_awaddr_s_o16                   =>  fabric_llpp3_awaddr_s_o(15)
       , fabric_llpp3_awaddr_s_o17                   =>  fabric_llpp3_awaddr_s_o(16)
       , fabric_llpp3_awaddr_s_o18                   =>  fabric_llpp3_awaddr_s_o(17)
       , fabric_llpp3_awaddr_s_o19                   =>  fabric_llpp3_awaddr_s_o(18)
       , fabric_llpp3_awaddr_s_o20                   =>  fabric_llpp3_awaddr_s_o(19)
       , fabric_llpp3_awaddr_s_o21                   =>  fabric_llpp3_awaddr_s_o(20)
       , fabric_llpp3_awaddr_s_o22                   =>  fabric_llpp3_awaddr_s_o(21)
       , fabric_llpp3_awaddr_s_o23                   =>  fabric_llpp3_awaddr_s_o(22)
       , fabric_llpp3_awaddr_s_o24                   =>  fabric_llpp3_awaddr_s_o(23)
       , fabric_llpp3_awaddr_s_o25                   =>  fabric_llpp3_awaddr_s_o(24)
       , fabric_llpp3_awaddr_s_o26                   =>  fabric_llpp3_awaddr_s_o(25)
       , fabric_llpp3_awaddr_s_o27                   =>  fabric_llpp3_awaddr_s_o(26)
       , fabric_llpp3_awaddr_s_o28                   =>  fabric_llpp3_awaddr_s_o(27)
       , fabric_llpp3_awaddr_s_o29                   =>  fabric_llpp3_awaddr_s_o(28)
       , fabric_llpp3_awaddr_s_o30                   =>  fabric_llpp3_awaddr_s_o(29)
       , fabric_llpp3_awaddr_s_o31                   =>  fabric_llpp3_awaddr_s_o(30)
       , fabric_llpp3_awaddr_s_o32                   =>  fabric_llpp3_awaddr_s_o(31)
       , fabric_llpp3_awburst_s_o1                   =>  fabric_llpp3_awburst_s_o(0)
       , fabric_llpp3_awburst_s_o2                   =>  fabric_llpp3_awburst_s_o(1)
       , fabric_llpp3_awcache_s_o1                   =>  fabric_llpp3_awcache_s_o(0)
       , fabric_llpp3_awcache_s_o2                   =>  fabric_llpp3_awcache_s_o(1)
       , fabric_llpp3_awcache_s_o3                   =>  fabric_llpp3_awcache_s_o(2)
       , fabric_llpp3_awcache_s_o4                   =>  fabric_llpp3_awcache_s_o(3)
       , fabric_llpp3_awid_s_o1                      =>  fabric_llpp3_awid_s_o(0)
       , fabric_llpp3_awid_s_o2                      =>  fabric_llpp3_awid_s_o(1)
       , fabric_llpp3_awid_s_o3                      =>  fabric_llpp3_awid_s_o(2)
       , fabric_llpp3_awid_s_o4                      =>  fabric_llpp3_awid_s_o(3)
       , fabric_llpp3_awid_s_o5                      =>  fabric_llpp3_awid_s_o(4)
       , fabric_llpp3_awid_s_o6                      =>  fabric_llpp3_awid_s_o(5)
       , fabric_llpp3_awid_s_o7                      =>  fabric_llpp3_awid_s_o(6)
       , fabric_llpp3_awid_s_o8                      =>  fabric_llpp3_awid_s_o(7)
       , fabric_llpp3_awid_s_o9                      =>  fabric_llpp3_awid_s_o(8)
       , fabric_llpp3_awid_s_o10                     =>  fabric_llpp3_awid_s_o(9)
       , fabric_llpp3_awid_s_o11                     =>  fabric_llpp3_awid_s_o(10)
       , fabric_llpp3_awid_s_o12                     =>  fabric_llpp3_awid_s_o(11)
       , fabric_llpp3_awlen_s_o1                     =>  fabric_llpp3_awlen_s_o(0)
       , fabric_llpp3_awlen_s_o2                     =>  fabric_llpp3_awlen_s_o(1)
       , fabric_llpp3_awlen_s_o3                     =>  fabric_llpp3_awlen_s_o(2)
       , fabric_llpp3_awlen_s_o4                     =>  fabric_llpp3_awlen_s_o(3)
       , fabric_llpp3_awlen_s_o5                     =>  fabric_llpp3_awlen_s_o(4)
       , fabric_llpp3_awlen_s_o6                     =>  fabric_llpp3_awlen_s_o(5)
       , fabric_llpp3_awlen_s_o7                     =>  fabric_llpp3_awlen_s_o(6)
       , fabric_llpp3_awlen_s_o8                     =>  fabric_llpp3_awlen_s_o(7)
       , fabric_llpp3_awlock_s_o                     =>  fabric_llpp3_awlock_s_o
       , fabric_llpp3_awprot_s_o1                    =>  fabric_llpp3_awprot_s_o(0)
       , fabric_llpp3_awprot_s_o2                    =>  fabric_llpp3_awprot_s_o(1)
       , fabric_llpp3_awprot_s_o3                    =>  fabric_llpp3_awprot_s_o(2)
       , fabric_llpp3_awqos_s_o1                     =>  fabric_llpp3_awqos_s_o(0)
       , fabric_llpp3_awqos_s_o2                     =>  fabric_llpp3_awqos_s_o(1)
       , fabric_llpp3_awqos_s_o3                     =>  fabric_llpp3_awqos_s_o(2)
       , fabric_llpp3_awqos_s_o4                     =>  fabric_llpp3_awqos_s_o(3)
       , fabric_llpp3_awsize_s_o1                    =>  fabric_llpp3_awsize_s_o(0)
       , fabric_llpp3_awsize_s_o2                    =>  fabric_llpp3_awsize_s_o(1)
       , fabric_llpp3_awsize_s_o3                    =>  fabric_llpp3_awsize_s_o(2)
       , fabric_llpp3_awvalid_s_o                    =>  fabric_llpp3_awvalid_s_o
       , fabric_llpp3_bready_s_o                     =>  fabric_llpp3_bready_s_o
       , fabric_llpp3_rready_s_o                     =>  fabric_llpp3_rready_s_o
       , fabric_llpp3_wdata_s_o1                     =>  fabric_llpp3_wdata_s_o(0)
       , fabric_llpp3_wdata_s_o2                     =>  fabric_llpp3_wdata_s_o(1)
       , fabric_llpp3_wdata_s_o3                     =>  fabric_llpp3_wdata_s_o(2)
       , fabric_llpp3_wdata_s_o4                     =>  fabric_llpp3_wdata_s_o(3)
       , fabric_llpp3_wdata_s_o5                     =>  fabric_llpp3_wdata_s_o(4)
       , fabric_llpp3_wdata_s_o6                     =>  fabric_llpp3_wdata_s_o(5)
       , fabric_llpp3_wdata_s_o7                     =>  fabric_llpp3_wdata_s_o(6)
       , fabric_llpp3_wdata_s_o8                     =>  fabric_llpp3_wdata_s_o(7)
       , fabric_llpp3_wdata_s_o9                     =>  fabric_llpp3_wdata_s_o(8)
       , fabric_llpp3_wdata_s_o10                    =>  fabric_llpp3_wdata_s_o(9)
       , fabric_llpp3_wdata_s_o11                    =>  fabric_llpp3_wdata_s_o(10)
       , fabric_llpp3_wdata_s_o12                    =>  fabric_llpp3_wdata_s_o(11)
       , fabric_llpp3_wdata_s_o13                    =>  fabric_llpp3_wdata_s_o(12)
       , fabric_llpp3_wdata_s_o14                    =>  fabric_llpp3_wdata_s_o(13)
       , fabric_llpp3_wdata_s_o15                    =>  fabric_llpp3_wdata_s_o(14)
       , fabric_llpp3_wdata_s_o16                    =>  fabric_llpp3_wdata_s_o(15)
       , fabric_llpp3_wdata_s_o17                    =>  fabric_llpp3_wdata_s_o(16)
       , fabric_llpp3_wdata_s_o18                    =>  fabric_llpp3_wdata_s_o(17)
       , fabric_llpp3_wdata_s_o19                    =>  fabric_llpp3_wdata_s_o(18)
       , fabric_llpp3_wdata_s_o20                    =>  fabric_llpp3_wdata_s_o(19)
       , fabric_llpp3_wdata_s_o21                    =>  fabric_llpp3_wdata_s_o(20)
       , fabric_llpp3_wdata_s_o22                    =>  fabric_llpp3_wdata_s_o(21)
       , fabric_llpp3_wdata_s_o23                    =>  fabric_llpp3_wdata_s_o(22)
       , fabric_llpp3_wdata_s_o24                    =>  fabric_llpp3_wdata_s_o(23)
       , fabric_llpp3_wdata_s_o25                    =>  fabric_llpp3_wdata_s_o(24)
       , fabric_llpp3_wdata_s_o26                    =>  fabric_llpp3_wdata_s_o(25)
       , fabric_llpp3_wdata_s_o27                    =>  fabric_llpp3_wdata_s_o(26)
       , fabric_llpp3_wdata_s_o28                    =>  fabric_llpp3_wdata_s_o(27)
       , fabric_llpp3_wdata_s_o29                    =>  fabric_llpp3_wdata_s_o(28)
       , fabric_llpp3_wdata_s_o30                    =>  fabric_llpp3_wdata_s_o(29)
       , fabric_llpp3_wdata_s_o31                    =>  fabric_llpp3_wdata_s_o(30)
       , fabric_llpp3_wdata_s_o32                    =>  fabric_llpp3_wdata_s_o(31)
       , fabric_llpp3_wlast_s_o                      =>  fabric_llpp3_wlast_s_o
       , fabric_llpp3_wstrb_s_o1                     =>  fabric_llpp3_wstrb_s_o(0)
       , fabric_llpp3_wstrb_s_o2                     =>  fabric_llpp3_wstrb_s_o(1)
       , fabric_llpp3_wstrb_s_o3                     =>  fabric_llpp3_wstrb_s_o(2)
       , fabric_llpp3_wstrb_s_o4                     =>  fabric_llpp3_wstrb_s_o(3)
       , fabric_llpp3_wvalid_s_o                     =>  fabric_llpp3_wvalid_s_o
       , fabric_llpp3_arready_s_i                    =>  fabric_llpp3_arready_s_i
       , fabric_llpp3_awready_s_i                    =>  fabric_llpp3_awready_s_i
       , fabric_llpp3_bid_s_i1                       =>  fabric_llpp3_bid_s_i(0)
       , fabric_llpp3_bid_s_i2                       =>  fabric_llpp3_bid_s_i(1)
       , fabric_llpp3_bid_s_i3                       =>  fabric_llpp3_bid_s_i(2)
       , fabric_llpp3_bid_s_i4                       =>  fabric_llpp3_bid_s_i(3)
       , fabric_llpp3_bid_s_i5                       =>  fabric_llpp3_bid_s_i(4)
       , fabric_llpp3_bid_s_i6                       =>  fabric_llpp3_bid_s_i(5)
       , fabric_llpp3_bid_s_i7                       =>  fabric_llpp3_bid_s_i(6)
       , fabric_llpp3_bid_s_i8                       =>  fabric_llpp3_bid_s_i(7)
       , fabric_llpp3_bid_s_i9                       =>  fabric_llpp3_bid_s_i(8)
       , fabric_llpp3_bid_s_i10                      =>  fabric_llpp3_bid_s_i(9)
       , fabric_llpp3_bid_s_i11                      =>  fabric_llpp3_bid_s_i(10)
       , fabric_llpp3_bid_s_i12                      =>  fabric_llpp3_bid_s_i(11)
       , fabric_llpp3_bresp_s_i1                     =>  fabric_llpp3_bresp_s_i(0)
       , fabric_llpp3_bresp_s_i2                     =>  fabric_llpp3_bresp_s_i(1)
       , fabric_llpp3_bvalid_s_i                     =>  fabric_llpp3_bvalid_s_i
       , fabric_llpp3_rdata_s_i1                     =>  fabric_llpp3_rdata_s_i(0)
       , fabric_llpp3_rdata_s_i2                     =>  fabric_llpp3_rdata_s_i(1)
       , fabric_llpp3_rdata_s_i3                     =>  fabric_llpp3_rdata_s_i(2)
       , fabric_llpp3_rdata_s_i4                     =>  fabric_llpp3_rdata_s_i(3)
       , fabric_llpp3_rdata_s_i5                     =>  fabric_llpp3_rdata_s_i(4)
       , fabric_llpp3_rdata_s_i6                     =>  fabric_llpp3_rdata_s_i(5)
       , fabric_llpp3_rdata_s_i7                     =>  fabric_llpp3_rdata_s_i(6)
       , fabric_llpp3_rdata_s_i8                     =>  fabric_llpp3_rdata_s_i(7)
       , fabric_llpp3_rdata_s_i9                     =>  fabric_llpp3_rdata_s_i(8)
       , fabric_llpp3_rdata_s_i10                    =>  fabric_llpp3_rdata_s_i(9)
       , fabric_llpp3_rdata_s_i11                    =>  fabric_llpp3_rdata_s_i(10)
       , fabric_llpp3_rdata_s_i12                    =>  fabric_llpp3_rdata_s_i(11)
       , fabric_llpp3_rdata_s_i13                    =>  fabric_llpp3_rdata_s_i(12)
       , fabric_llpp3_rdata_s_i14                    =>  fabric_llpp3_rdata_s_i(13)
       , fabric_llpp3_rdata_s_i15                    =>  fabric_llpp3_rdata_s_i(14)
       , fabric_llpp3_rdata_s_i16                    =>  fabric_llpp3_rdata_s_i(15)
       , fabric_llpp3_rdata_s_i17                    =>  fabric_llpp3_rdata_s_i(16)
       , fabric_llpp3_rdata_s_i18                    =>  fabric_llpp3_rdata_s_i(17)
       , fabric_llpp3_rdata_s_i19                    =>  fabric_llpp3_rdata_s_i(18)
       , fabric_llpp3_rdata_s_i20                    =>  fabric_llpp3_rdata_s_i(19)
       , fabric_llpp3_rdata_s_i21                    =>  fabric_llpp3_rdata_s_i(20)
       , fabric_llpp3_rdata_s_i22                    =>  fabric_llpp3_rdata_s_i(21)
       , fabric_llpp3_rdata_s_i23                    =>  fabric_llpp3_rdata_s_i(22)
       , fabric_llpp3_rdata_s_i24                    =>  fabric_llpp3_rdata_s_i(23)
       , fabric_llpp3_rdata_s_i25                    =>  fabric_llpp3_rdata_s_i(24)
       , fabric_llpp3_rdata_s_i26                    =>  fabric_llpp3_rdata_s_i(25)
       , fabric_llpp3_rdata_s_i27                    =>  fabric_llpp3_rdata_s_i(26)
       , fabric_llpp3_rdata_s_i28                    =>  fabric_llpp3_rdata_s_i(27)
       , fabric_llpp3_rdata_s_i29                    =>  fabric_llpp3_rdata_s_i(28)
       , fabric_llpp3_rdata_s_i30                    =>  fabric_llpp3_rdata_s_i(29)
       , fabric_llpp3_rdata_s_i31                    =>  fabric_llpp3_rdata_s_i(30)
       , fabric_llpp3_rdata_s_i32                    =>  fabric_llpp3_rdata_s_i(31)
       , fabric_llpp3_rid_s_i1                       =>  fabric_llpp3_rid_s_i(0)
       , fabric_llpp3_rid_s_i2                       =>  fabric_llpp3_rid_s_i(1)
       , fabric_llpp3_rid_s_i3                       =>  fabric_llpp3_rid_s_i(2)
       , fabric_llpp3_rid_s_i4                       =>  fabric_llpp3_rid_s_i(3)
       , fabric_llpp3_rid_s_i5                       =>  fabric_llpp3_rid_s_i(4)
       , fabric_llpp3_rid_s_i6                       =>  fabric_llpp3_rid_s_i(5)
       , fabric_llpp3_rid_s_i7                       =>  fabric_llpp3_rid_s_i(6)
       , fabric_llpp3_rid_s_i8                       =>  fabric_llpp3_rid_s_i(7)
       , fabric_llpp3_rid_s_i9                       =>  fabric_llpp3_rid_s_i(8)
       , fabric_llpp3_rid_s_i10                      =>  fabric_llpp3_rid_s_i(9)
       , fabric_llpp3_rid_s_i11                      =>  fabric_llpp3_rid_s_i(10)
       , fabric_llpp3_rid_s_i12                      =>  fabric_llpp3_rid_s_i(11)
       , fabric_llpp3_rlast_s_i                      =>  fabric_llpp3_rlast_s_i
       , fabric_llpp3_rresp_s_i1                     =>  fabric_llpp3_rresp_s_i(0)
       , fabric_llpp3_rresp_s_i2                     =>  fabric_llpp3_rresp_s_i(1)
       , fabric_llpp3_rvalid_s_i                     =>  fabric_llpp3_rvalid_s_i
       , fabric_llpp3_wready_s_i                     =>  fabric_llpp3_wready_s_i
       , fabric_qos_pprdata_o1                       =>  fabric_qos_pprdata_o(0)
       , fabric_qos_pprdata_o2                       =>  fabric_qos_pprdata_o(1)
       , fabric_qos_pprdata_o3                       =>  fabric_qos_pprdata_o(2)
       , fabric_qos_pprdata_o4                       =>  fabric_qos_pprdata_o(3)
       , fabric_qos_pprdata_o5                       =>  fabric_qos_pprdata_o(4)
       , fabric_qos_pprdata_o6                       =>  fabric_qos_pprdata_o(5)
       , fabric_qos_pprdata_o7                       =>  fabric_qos_pprdata_o(6)
       , fabric_qos_pprdata_o8                       =>  fabric_qos_pprdata_o(7)
       , fabric_qos_pprdata_o9                       =>  fabric_qos_pprdata_o(8)
       , fabric_qos_pprdata_o10                      =>  fabric_qos_pprdata_o(9)
       , fabric_qos_pprdata_o11                      =>  fabric_qos_pprdata_o(10)
       , fabric_qos_pprdata_o12                      =>  fabric_qos_pprdata_o(11)
       , fabric_qos_pprdata_o13                      =>  fabric_qos_pprdata_o(12)
       , fabric_qos_pprdata_o14                      =>  fabric_qos_pprdata_o(13)
       , fabric_qos_pprdata_o15                      =>  fabric_qos_pprdata_o(14)
       , fabric_qos_pprdata_o16                      =>  fabric_qos_pprdata_o(15)
       , fabric_qos_pprdata_o17                      =>  fabric_qos_pprdata_o(16)
       , fabric_qos_pprdata_o18                      =>  fabric_qos_pprdata_o(17)
       , fabric_qos_pprdata_o19                      =>  fabric_qos_pprdata_o(18)
       , fabric_qos_pprdata_o20                      =>  fabric_qos_pprdata_o(19)
       , fabric_qos_pprdata_o21                      =>  fabric_qos_pprdata_o(20)
       , fabric_qos_pprdata_o22                      =>  fabric_qos_pprdata_o(21)
       , fabric_qos_pprdata_o23                      =>  fabric_qos_pprdata_o(22)
       , fabric_qos_pprdata_o24                      =>  fabric_qos_pprdata_o(23)
       , fabric_qos_pprdata_o25                      =>  fabric_qos_pprdata_o(24)
       , fabric_qos_pprdata_o26                      =>  fabric_qos_pprdata_o(25)
       , fabric_qos_pprdata_o27                      =>  fabric_qos_pprdata_o(26)
       , fabric_qos_pprdata_o28                      =>  fabric_qos_pprdata_o(27)
       , fabric_qos_pprdata_o29                      =>  fabric_qos_pprdata_o(28)
       , fabric_qos_pprdata_o30                      =>  fabric_qos_pprdata_o(29)
       , fabric_qos_pprdata_o31                      =>  fabric_qos_pprdata_o(30)
       , fabric_qos_pprdata_o32                      =>  fabric_qos_pprdata_o(31)
       , fabric_qos_ppready_o                        =>  fabric_qos_ppready_o
       , fabric_qos_ppslverr_o                       =>  fabric_qos_ppslverr_o
       , fabric_qos_pclk_i                           =>  fabric_qos_pclk_i
       , fabric_qos_ppaddr_i1                        =>  fabric_qos_ppaddr_i(0)
       , fabric_qos_ppaddr_i2                        =>  fabric_qos_ppaddr_i(1)
       , fabric_qos_ppaddr_i3                        =>  fabric_qos_ppaddr_i(2)
       , fabric_qos_ppaddr_i4                        =>  fabric_qos_ppaddr_i(3)
       , fabric_qos_ppaddr_i5                        =>  fabric_qos_ppaddr_i(4)
       , fabric_qos_ppaddr_i6                        =>  fabric_qos_ppaddr_i(5)
       , fabric_qos_ppaddr_i7                        =>  fabric_qos_ppaddr_i(6)
       , fabric_qos_ppaddr_i8                        =>  fabric_qos_ppaddr_i(7)
       , fabric_qos_ppaddr_i9                        =>  fabric_qos_ppaddr_i(8)
       , fabric_qos_ppaddr_i10                       =>  fabric_qos_ppaddr_i(9)
       , fabric_qos_ppaddr_i11                       =>  fabric_qos_ppaddr_i(10)
       , fabric_qos_ppaddr_i12                       =>  fabric_qos_ppaddr_i(11)
       , fabric_qos_ppaddr_i13                       =>  fabric_qos_ppaddr_i(12)
       , fabric_qos_ppaddr_i14                       =>  fabric_qos_ppaddr_i(13)
       , fabric_qos_ppaddr_i15                       =>  fabric_qos_ppaddr_i(14)
       , fabric_qos_ppaddr_i16                       =>  fabric_qos_ppaddr_i(15)
       , fabric_qos_ppaddr_i17                       =>  fabric_qos_ppaddr_i(16)
       , fabric_qos_ppaddr_i18                       =>  fabric_qos_ppaddr_i(17)
       , fabric_qos_ppaddr_i19                       =>  fabric_qos_ppaddr_i(18)
       , fabric_qos_ppaddr_i20                       =>  fabric_qos_ppaddr_i(19)
       , fabric_qos_ppaddr_i21                       =>  fabric_qos_ppaddr_i(20)
       , fabric_qos_ppaddr_i22                       =>  fabric_qos_ppaddr_i(21)
       , fabric_qos_ppaddr_i23                       =>  fabric_qos_ppaddr_i(22)
       , fabric_qos_ppaddr_i24                       =>  fabric_qos_ppaddr_i(23)
       , fabric_qos_ppaddr_i25                       =>  fabric_qos_ppaddr_i(24)
       , fabric_qos_ppaddr_i26                       =>  fabric_qos_ppaddr_i(25)
       , fabric_qos_ppaddr_i27                       =>  fabric_qos_ppaddr_i(26)
       , fabric_qos_ppaddr_i28                       =>  fabric_qos_ppaddr_i(27)
       , fabric_qos_ppaddr_i29                       =>  fabric_qos_ppaddr_i(28)
       , fabric_qos_ppaddr_i30                       =>  fabric_qos_ppaddr_i(29)
       , fabric_qos_ppaddr_i31                       =>  fabric_qos_ppaddr_i(30)
       , fabric_qos_ppaddr_i32                       =>  fabric_qos_ppaddr_i(31)
       , fabric_qos_ppenable_i                       =>  fabric_qos_ppenable_i
       , fabric_qos_ppwdata_i1                       =>  fabric_qos_ppwdata_i(0)
       , fabric_qos_ppwdata_i2                       =>  fabric_qos_ppwdata_i(1)
       , fabric_qos_ppwdata_i3                       =>  fabric_qos_ppwdata_i(2)
       , fabric_qos_ppwdata_i4                       =>  fabric_qos_ppwdata_i(3)
       , fabric_qos_ppwdata_i5                       =>  fabric_qos_ppwdata_i(4)
       , fabric_qos_ppwdata_i6                       =>  fabric_qos_ppwdata_i(5)
       , fabric_qos_ppwdata_i7                       =>  fabric_qos_ppwdata_i(6)
       , fabric_qos_ppwdata_i8                       =>  fabric_qos_ppwdata_i(7)
       , fabric_qos_ppwdata_i9                       =>  fabric_qos_ppwdata_i(8)
       , fabric_qos_ppwdata_i10                      =>  fabric_qos_ppwdata_i(9)
       , fabric_qos_ppwdata_i11                      =>  fabric_qos_ppwdata_i(10)
       , fabric_qos_ppwdata_i12                      =>  fabric_qos_ppwdata_i(11)
       , fabric_qos_ppwdata_i13                      =>  fabric_qos_ppwdata_i(12)
       , fabric_qos_ppwdata_i14                      =>  fabric_qos_ppwdata_i(13)
       , fabric_qos_ppwdata_i15                      =>  fabric_qos_ppwdata_i(14)
       , fabric_qos_ppwdata_i16                      =>  fabric_qos_ppwdata_i(15)
       , fabric_qos_ppwdata_i17                      =>  fabric_qos_ppwdata_i(16)
       , fabric_qos_ppwdata_i18                      =>  fabric_qos_ppwdata_i(17)
       , fabric_qos_ppwdata_i19                      =>  fabric_qos_ppwdata_i(18)
       , fabric_qos_ppwdata_i20                      =>  fabric_qos_ppwdata_i(19)
       , fabric_qos_ppwdata_i21                      =>  fabric_qos_ppwdata_i(20)
       , fabric_qos_ppwdata_i22                      =>  fabric_qos_ppwdata_i(21)
       , fabric_qos_ppwdata_i23                      =>  fabric_qos_ppwdata_i(22)
       , fabric_qos_ppwdata_i24                      =>  fabric_qos_ppwdata_i(23)
       , fabric_qos_ppwdata_i25                      =>  fabric_qos_ppwdata_i(24)
       , fabric_qos_ppwdata_i26                      =>  fabric_qos_ppwdata_i(25)
       , fabric_qos_ppwdata_i27                      =>  fabric_qos_ppwdata_i(26)
       , fabric_qos_ppwdata_i28                      =>  fabric_qos_ppwdata_i(27)
       , fabric_qos_ppwdata_i29                      =>  fabric_qos_ppwdata_i(28)
       , fabric_qos_ppwdata_i30                      =>  fabric_qos_ppwdata_i(29)
       , fabric_qos_ppwdata_i31                      =>  fabric_qos_ppwdata_i(30)
       , fabric_qos_ppwdata_i32                      =>  fabric_qos_ppwdata_i(31)
       , fabric_qos_ppwrite_i                        =>  fabric_qos_ppwrite_i
       , fabric_qos_presetn_i                        =>  fabric_qos_presetn_i
       , fabric_qos_psel_i                           =>  fabric_qos_psel_i
       , fabric_tnd_hssl_flushin_o                   =>  fabric_tnd_hssl_flushin_o
       , fabric_tnd_hssl_trigin_o                    =>  fabric_tnd_hssl_trigin_o
       , fabric_tnd_fpga_apb_master_paddr_o1         =>  fabric_tnd_fpga_apb_master_paddr_o(0)
       , fabric_tnd_fpga_apb_master_paddr_o2         =>  fabric_tnd_fpga_apb_master_paddr_o(1)
       , fabric_tnd_fpga_apb_master_paddr_o3         =>  fabric_tnd_fpga_apb_master_paddr_o(2)
       , fabric_tnd_fpga_apb_master_paddr_o4         =>  fabric_tnd_fpga_apb_master_paddr_o(3)
       , fabric_tnd_fpga_apb_master_paddr_o5         =>  fabric_tnd_fpga_apb_master_paddr_o(4)
       , fabric_tnd_fpga_apb_master_paddr_o6         =>  fabric_tnd_fpga_apb_master_paddr_o(5)
       , fabric_tnd_fpga_apb_master_paddr_o7         =>  fabric_tnd_fpga_apb_master_paddr_o(6)
       , fabric_tnd_fpga_apb_master_paddr_o8         =>  fabric_tnd_fpga_apb_master_paddr_o(7)
       , fabric_tnd_fpga_apb_master_paddr_o9         =>  fabric_tnd_fpga_apb_master_paddr_o(8)
       , fabric_tnd_fpga_apb_master_paddr_o10        =>  fabric_tnd_fpga_apb_master_paddr_o(9)
       , fabric_tnd_fpga_apb_master_paddr_o11        =>  fabric_tnd_fpga_apb_master_paddr_o(10)
       , fabric_tnd_fpga_apb_master_paddr_o12        =>  fabric_tnd_fpga_apb_master_paddr_o(11)
       , fabric_tnd_fpga_apb_master_paddr_o13        =>  fabric_tnd_fpga_apb_master_paddr_o(12)
       , fabric_tnd_fpga_apb_master_paddr_o14        =>  fabric_tnd_fpga_apb_master_paddr_o(13)
       , fabric_tnd_fpga_apb_master_paddr_o15        =>  fabric_tnd_fpga_apb_master_paddr_o(14)
       , fabric_tnd_fpga_apb_master_paddr_o16        =>  fabric_tnd_fpga_apb_master_paddr_o(15)
       , fabric_tnd_fpga_apb_master_paddr_o17        =>  fabric_tnd_fpga_apb_master_paddr_o(16)
       , fabric_tnd_fpga_apb_master_paddr_o18        =>  fabric_tnd_fpga_apb_master_paddr_o(17)
       , fabric_tnd_fpga_apb_master_paddr_o19        =>  fabric_tnd_fpga_apb_master_paddr_o(18)
       , fabric_tnd_fpga_apb_master_paddr_o20        =>  fabric_tnd_fpga_apb_master_paddr_o(19)
       , fabric_tnd_fpga_apb_master_paddr_o21        =>  fabric_tnd_fpga_apb_master_paddr_o(20)
       , fabric_tnd_fpga_apb_master_paddr_o22        =>  fabric_tnd_fpga_apb_master_paddr_o(21)
       , fabric_tnd_fpga_apb_master_paddr_o23        =>  fabric_tnd_fpga_apb_master_paddr_o(22)
       , fabric_tnd_fpga_apb_master_paddr_o24        =>  fabric_tnd_fpga_apb_master_paddr_o(23)
       , fabric_tnd_fpga_apb_master_paddr_o25        =>  fabric_tnd_fpga_apb_master_paddr_o(24)
       , fabric_tnd_fpga_apb_master_paddr_o26        =>  fabric_tnd_fpga_apb_master_paddr_o(25)
       , fabric_tnd_fpga_apb_master_paddr_o27        =>  fabric_tnd_fpga_apb_master_paddr_o(26)
       , fabric_tnd_fpga_apb_master_paddr_o28        =>  fabric_tnd_fpga_apb_master_paddr_o(27)
       , fabric_tnd_fpga_apb_master_paddr_o29        =>  fabric_tnd_fpga_apb_master_paddr_o(28)
       , fabric_tnd_fpga_apb_master_paddr_o30        =>  fabric_tnd_fpga_apb_master_paddr_o(29)
       , fabric_tnd_fpga_apb_master_paddr_o31        =>  fabric_tnd_fpga_apb_master_paddr_o(30)
       , fabric_tnd_fpga_apb_master_paddr_o32        =>  fabric_tnd_fpga_apb_master_paddr_o(31)
       , fabric_tnd_fpga_apb_master_penable_o        =>  fabric_tnd_fpga_apb_master_penable_o
       , fabric_tnd_fpga_apb_master_psel_o           =>  fabric_tnd_fpga_apb_master_psel_o
       , fabric_tnd_fpga_apb_master_pwdata_o1        =>  fabric_tnd_fpga_apb_master_pwdata_o(0)
       , fabric_tnd_fpga_apb_master_pwdata_o2        =>  fabric_tnd_fpga_apb_master_pwdata_o(1)
       , fabric_tnd_fpga_apb_master_pwdata_o3        =>  fabric_tnd_fpga_apb_master_pwdata_o(2)
       , fabric_tnd_fpga_apb_master_pwdata_o4        =>  fabric_tnd_fpga_apb_master_pwdata_o(3)
       , fabric_tnd_fpga_apb_master_pwdata_o5        =>  fabric_tnd_fpga_apb_master_pwdata_o(4)
       , fabric_tnd_fpga_apb_master_pwdata_o6        =>  fabric_tnd_fpga_apb_master_pwdata_o(5)
       , fabric_tnd_fpga_apb_master_pwdata_o7        =>  fabric_tnd_fpga_apb_master_pwdata_o(6)
       , fabric_tnd_fpga_apb_master_pwdata_o8        =>  fabric_tnd_fpga_apb_master_pwdata_o(7)
       , fabric_tnd_fpga_apb_master_pwdata_o9        =>  fabric_tnd_fpga_apb_master_pwdata_o(8)
       , fabric_tnd_fpga_apb_master_pwdata_o10       =>  fabric_tnd_fpga_apb_master_pwdata_o(9)
       , fabric_tnd_fpga_apb_master_pwdata_o11       =>  fabric_tnd_fpga_apb_master_pwdata_o(10)
       , fabric_tnd_fpga_apb_master_pwdata_o12       =>  fabric_tnd_fpga_apb_master_pwdata_o(11)
       , fabric_tnd_fpga_apb_master_pwdata_o13       =>  fabric_tnd_fpga_apb_master_pwdata_o(12)
       , fabric_tnd_fpga_apb_master_pwdata_o14       =>  fabric_tnd_fpga_apb_master_pwdata_o(13)
       , fabric_tnd_fpga_apb_master_pwdata_o15       =>  fabric_tnd_fpga_apb_master_pwdata_o(14)
       , fabric_tnd_fpga_apb_master_pwdata_o16       =>  fabric_tnd_fpga_apb_master_pwdata_o(15)
       , fabric_tnd_fpga_apb_master_pwdata_o17       =>  fabric_tnd_fpga_apb_master_pwdata_o(16)
       , fabric_tnd_fpga_apb_master_pwdata_o18       =>  fabric_tnd_fpga_apb_master_pwdata_o(17)
       , fabric_tnd_fpga_apb_master_pwdata_o19       =>  fabric_tnd_fpga_apb_master_pwdata_o(18)
       , fabric_tnd_fpga_apb_master_pwdata_o20       =>  fabric_tnd_fpga_apb_master_pwdata_o(19)
       , fabric_tnd_fpga_apb_master_pwdata_o21       =>  fabric_tnd_fpga_apb_master_pwdata_o(20)
       , fabric_tnd_fpga_apb_master_pwdata_o22       =>  fabric_tnd_fpga_apb_master_pwdata_o(21)
       , fabric_tnd_fpga_apb_master_pwdata_o23       =>  fabric_tnd_fpga_apb_master_pwdata_o(22)
       , fabric_tnd_fpga_apb_master_pwdata_o24       =>  fabric_tnd_fpga_apb_master_pwdata_o(23)
       , fabric_tnd_fpga_apb_master_pwdata_o25       =>  fabric_tnd_fpga_apb_master_pwdata_o(24)
       , fabric_tnd_fpga_apb_master_pwdata_o26       =>  fabric_tnd_fpga_apb_master_pwdata_o(25)
       , fabric_tnd_fpga_apb_master_pwdata_o27       =>  fabric_tnd_fpga_apb_master_pwdata_o(26)
       , fabric_tnd_fpga_apb_master_pwdata_o28       =>  fabric_tnd_fpga_apb_master_pwdata_o(27)
       , fabric_tnd_fpga_apb_master_pwdata_o29       =>  fabric_tnd_fpga_apb_master_pwdata_o(28)
       , fabric_tnd_fpga_apb_master_pwdata_o30       =>  fabric_tnd_fpga_apb_master_pwdata_o(29)
       , fabric_tnd_fpga_apb_master_pwdata_o31       =>  fabric_tnd_fpga_apb_master_pwdata_o(30)
       , fabric_tnd_fpga_apb_master_pwdata_o32       =>  fabric_tnd_fpga_apb_master_pwdata_o(31)
       , fabric_tnd_fpga_apb_master_pwrite_o         =>  fabric_tnd_fpga_apb_master_pwrite_o
       , fabric_tnd_fpga_atb_master_afvalid_o        =>  fabric_tnd_fpga_atb_master_afvalid_o
       , fabric_tnd_fpga_atb_master_atready_o        =>  fabric_tnd_fpga_atb_master_atready_o
       , fabric_tnd_fpga_atb_master_syncreq_o        =>  fabric_tnd_fpga_atb_master_syncreq_o
       , fabric_tnd_hssl_apb_master_paddr_o1         =>  fabric_tnd_hssl_apb_master_paddr_o(0)
       , fabric_tnd_hssl_apb_master_paddr_o2         =>  fabric_tnd_hssl_apb_master_paddr_o(1)
       , fabric_tnd_hssl_apb_master_paddr_o3         =>  fabric_tnd_hssl_apb_master_paddr_o(2)
       , fabric_tnd_hssl_apb_master_paddr_o4         =>  fabric_tnd_hssl_apb_master_paddr_o(3)
       , fabric_tnd_hssl_apb_master_paddr_o5         =>  fabric_tnd_hssl_apb_master_paddr_o(4)
       , fabric_tnd_hssl_apb_master_paddr_o6         =>  fabric_tnd_hssl_apb_master_paddr_o(5)
       , fabric_tnd_hssl_apb_master_paddr_o7         =>  fabric_tnd_hssl_apb_master_paddr_o(6)
       , fabric_tnd_hssl_apb_master_paddr_o8         =>  fabric_tnd_hssl_apb_master_paddr_o(7)
       , fabric_tnd_hssl_apb_master_paddr_o9         =>  fabric_tnd_hssl_apb_master_paddr_o(8)
       , fabric_tnd_hssl_apb_master_paddr_o10        =>  fabric_tnd_hssl_apb_master_paddr_o(9)
       , fabric_tnd_hssl_apb_master_paddr_o11        =>  fabric_tnd_hssl_apb_master_paddr_o(10)
       , fabric_tnd_hssl_apb_master_paddr_o12        =>  fabric_tnd_hssl_apb_master_paddr_o(11)
       , fabric_tnd_hssl_apb_master_paddr_o13        =>  fabric_tnd_hssl_apb_master_paddr_o(12)
       , fabric_tnd_hssl_apb_master_paddr_o14        =>  fabric_tnd_hssl_apb_master_paddr_o(13)
       , fabric_tnd_hssl_apb_master_paddr_o15        =>  fabric_tnd_hssl_apb_master_paddr_o(14)
       , fabric_tnd_hssl_apb_master_paddr_o16        =>  fabric_tnd_hssl_apb_master_paddr_o(15)
       , fabric_tnd_hssl_apb_master_paddr_o17        =>  fabric_tnd_hssl_apb_master_paddr_o(16)
       , fabric_tnd_hssl_apb_master_paddr_o18        =>  fabric_tnd_hssl_apb_master_paddr_o(17)
       , fabric_tnd_hssl_apb_master_paddr_o19        =>  fabric_tnd_hssl_apb_master_paddr_o(18)
       , fabric_tnd_hssl_apb_master_paddr_o20        =>  fabric_tnd_hssl_apb_master_paddr_o(19)
       , fabric_tnd_hssl_apb_master_paddr_o21        =>  fabric_tnd_hssl_apb_master_paddr_o(20)
       , fabric_tnd_hssl_apb_master_paddr_o22        =>  fabric_tnd_hssl_apb_master_paddr_o(21)
       , fabric_tnd_hssl_apb_master_paddr_o23        =>  fabric_tnd_hssl_apb_master_paddr_o(22)
       , fabric_tnd_hssl_apb_master_paddr_o24        =>  fabric_tnd_hssl_apb_master_paddr_o(23)
       , fabric_tnd_hssl_apb_master_paddr_o25        =>  fabric_tnd_hssl_apb_master_paddr_o(24)
       , fabric_tnd_hssl_apb_master_paddr_o26        =>  fabric_tnd_hssl_apb_master_paddr_o(25)
       , fabric_tnd_hssl_apb_master_paddr_o27        =>  fabric_tnd_hssl_apb_master_paddr_o(26)
       , fabric_tnd_hssl_apb_master_paddr_o28        =>  fabric_tnd_hssl_apb_master_paddr_o(27)
       , fabric_tnd_hssl_apb_master_paddr_o29        =>  fabric_tnd_hssl_apb_master_paddr_o(28)
       , fabric_tnd_hssl_apb_master_paddr_o30        =>  fabric_tnd_hssl_apb_master_paddr_o(29)
       , fabric_tnd_hssl_apb_master_paddr_o31        =>  fabric_tnd_hssl_apb_master_paddr_o(30)
       , fabric_tnd_hssl_apb_master_paddr_o32        =>  fabric_tnd_hssl_apb_master_paddr_o(31)
       , fabric_tnd_hssl_apb_master_penable_o        =>  fabric_tnd_hssl_apb_master_penable_o
       , fabric_tnd_hssl_apb_master_psel_o           =>  fabric_tnd_hssl_apb_master_psel_o
       , fabric_tnd_hssl_apb_master_pwdata_o1        =>  fabric_tnd_hssl_apb_master_pwdata_o(0)
       , fabric_tnd_hssl_apb_master_pwdata_o2        =>  fabric_tnd_hssl_apb_master_pwdata_o(1)
       , fabric_tnd_hssl_apb_master_pwdata_o3        =>  fabric_tnd_hssl_apb_master_pwdata_o(2)
       , fabric_tnd_hssl_apb_master_pwdata_o4        =>  fabric_tnd_hssl_apb_master_pwdata_o(3)
       , fabric_tnd_hssl_apb_master_pwdata_o5        =>  fabric_tnd_hssl_apb_master_pwdata_o(4)
       , fabric_tnd_hssl_apb_master_pwdata_o6        =>  fabric_tnd_hssl_apb_master_pwdata_o(5)
       , fabric_tnd_hssl_apb_master_pwdata_o7        =>  fabric_tnd_hssl_apb_master_pwdata_o(6)
       , fabric_tnd_hssl_apb_master_pwdata_o8        =>  fabric_tnd_hssl_apb_master_pwdata_o(7)
       , fabric_tnd_hssl_apb_master_pwdata_o9        =>  fabric_tnd_hssl_apb_master_pwdata_o(8)
       , fabric_tnd_hssl_apb_master_pwdata_o10       =>  fabric_tnd_hssl_apb_master_pwdata_o(9)
       , fabric_tnd_hssl_apb_master_pwdata_o11       =>  fabric_tnd_hssl_apb_master_pwdata_o(10)
       , fabric_tnd_hssl_apb_master_pwdata_o12       =>  fabric_tnd_hssl_apb_master_pwdata_o(11)
       , fabric_tnd_hssl_apb_master_pwdata_o13       =>  fabric_tnd_hssl_apb_master_pwdata_o(12)
       , fabric_tnd_hssl_apb_master_pwdata_o14       =>  fabric_tnd_hssl_apb_master_pwdata_o(13)
       , fabric_tnd_hssl_apb_master_pwdata_o15       =>  fabric_tnd_hssl_apb_master_pwdata_o(14)
       , fabric_tnd_hssl_apb_master_pwdata_o16       =>  fabric_tnd_hssl_apb_master_pwdata_o(15)
       , fabric_tnd_hssl_apb_master_pwdata_o17       =>  fabric_tnd_hssl_apb_master_pwdata_o(16)
       , fabric_tnd_hssl_apb_master_pwdata_o18       =>  fabric_tnd_hssl_apb_master_pwdata_o(17)
       , fabric_tnd_hssl_apb_master_pwdata_o19       =>  fabric_tnd_hssl_apb_master_pwdata_o(18)
       , fabric_tnd_hssl_apb_master_pwdata_o20       =>  fabric_tnd_hssl_apb_master_pwdata_o(19)
       , fabric_tnd_hssl_apb_master_pwdata_o21       =>  fabric_tnd_hssl_apb_master_pwdata_o(20)
       , fabric_tnd_hssl_apb_master_pwdata_o22       =>  fabric_tnd_hssl_apb_master_pwdata_o(21)
       , fabric_tnd_hssl_apb_master_pwdata_o23       =>  fabric_tnd_hssl_apb_master_pwdata_o(22)
       , fabric_tnd_hssl_apb_master_pwdata_o24       =>  fabric_tnd_hssl_apb_master_pwdata_o(23)
       , fabric_tnd_hssl_apb_master_pwdata_o25       =>  fabric_tnd_hssl_apb_master_pwdata_o(24)
       , fabric_tnd_hssl_apb_master_pwdata_o26       =>  fabric_tnd_hssl_apb_master_pwdata_o(25)
       , fabric_tnd_hssl_apb_master_pwdata_o27       =>  fabric_tnd_hssl_apb_master_pwdata_o(26)
       , fabric_tnd_hssl_apb_master_pwdata_o28       =>  fabric_tnd_hssl_apb_master_pwdata_o(27)
       , fabric_tnd_hssl_apb_master_pwdata_o29       =>  fabric_tnd_hssl_apb_master_pwdata_o(28)
       , fabric_tnd_hssl_apb_master_pwdata_o30       =>  fabric_tnd_hssl_apb_master_pwdata_o(29)
       , fabric_tnd_hssl_apb_master_pwdata_o31       =>  fabric_tnd_hssl_apb_master_pwdata_o(30)
       , fabric_tnd_hssl_apb_master_pwdata_o32       =>  fabric_tnd_hssl_apb_master_pwdata_o(31)
       , fabric_tnd_hssl_apb_master_pwrite_o         =>  fabric_tnd_hssl_apb_master_pwrite_o
       , fabric_tnd_hssl_atb_master_afready_o        =>  fabric_tnd_hssl_atb_master_afready_o
       , fabric_tnd_hssl_atb_master_atbytes_o1       =>  fabric_tnd_hssl_atb_master_atbytes_o(0)
       , fabric_tnd_hssl_atb_master_atbytes_o2       =>  fabric_tnd_hssl_atb_master_atbytes_o(1)
       , fabric_tnd_hssl_atb_master_atbytes_o3       =>  fabric_tnd_hssl_atb_master_atbytes_o(2)
       , fabric_tnd_hssl_atb_master_atbytes_o4       =>  fabric_tnd_hssl_atb_master_atbytes_o(3)
       , fabric_tnd_hssl_atb_master_atdata_o1        =>  fabric_tnd_hssl_atb_master_atdata_o(0)
       , fabric_tnd_hssl_atb_master_atdata_o2        =>  fabric_tnd_hssl_atb_master_atdata_o(1)
       , fabric_tnd_hssl_atb_master_atdata_o3        =>  fabric_tnd_hssl_atb_master_atdata_o(2)
       , fabric_tnd_hssl_atb_master_atdata_o4        =>  fabric_tnd_hssl_atb_master_atdata_o(3)
       , fabric_tnd_hssl_atb_master_atdata_o5        =>  fabric_tnd_hssl_atb_master_atdata_o(4)
       , fabric_tnd_hssl_atb_master_atdata_o6        =>  fabric_tnd_hssl_atb_master_atdata_o(5)
       , fabric_tnd_hssl_atb_master_atdata_o7        =>  fabric_tnd_hssl_atb_master_atdata_o(6)
       , fabric_tnd_hssl_atb_master_atdata_o8        =>  fabric_tnd_hssl_atb_master_atdata_o(7)
       , fabric_tnd_hssl_atb_master_atdata_o9        =>  fabric_tnd_hssl_atb_master_atdata_o(8)
       , fabric_tnd_hssl_atb_master_atdata_o10       =>  fabric_tnd_hssl_atb_master_atdata_o(9)
       , fabric_tnd_hssl_atb_master_atdata_o11       =>  fabric_tnd_hssl_atb_master_atdata_o(10)
       , fabric_tnd_hssl_atb_master_atdata_o12       =>  fabric_tnd_hssl_atb_master_atdata_o(11)
       , fabric_tnd_hssl_atb_master_atdata_o13       =>  fabric_tnd_hssl_atb_master_atdata_o(12)
       , fabric_tnd_hssl_atb_master_atdata_o14       =>  fabric_tnd_hssl_atb_master_atdata_o(13)
       , fabric_tnd_hssl_atb_master_atdata_o15       =>  fabric_tnd_hssl_atb_master_atdata_o(14)
       , fabric_tnd_hssl_atb_master_atdata_o16       =>  fabric_tnd_hssl_atb_master_atdata_o(15)
       , fabric_tnd_hssl_atb_master_atdata_o17       =>  fabric_tnd_hssl_atb_master_atdata_o(16)
       , fabric_tnd_hssl_atb_master_atdata_o18       =>  fabric_tnd_hssl_atb_master_atdata_o(17)
       , fabric_tnd_hssl_atb_master_atdata_o19       =>  fabric_tnd_hssl_atb_master_atdata_o(18)
       , fabric_tnd_hssl_atb_master_atdata_o20       =>  fabric_tnd_hssl_atb_master_atdata_o(19)
       , fabric_tnd_hssl_atb_master_atdata_o21       =>  fabric_tnd_hssl_atb_master_atdata_o(20)
       , fabric_tnd_hssl_atb_master_atdata_o22       =>  fabric_tnd_hssl_atb_master_atdata_o(21)
       , fabric_tnd_hssl_atb_master_atdata_o23       =>  fabric_tnd_hssl_atb_master_atdata_o(22)
       , fabric_tnd_hssl_atb_master_atdata_o24       =>  fabric_tnd_hssl_atb_master_atdata_o(23)
       , fabric_tnd_hssl_atb_master_atdata_o25       =>  fabric_tnd_hssl_atb_master_atdata_o(24)
       , fabric_tnd_hssl_atb_master_atdata_o26       =>  fabric_tnd_hssl_atb_master_atdata_o(25)
       , fabric_tnd_hssl_atb_master_atdata_o27       =>  fabric_tnd_hssl_atb_master_atdata_o(26)
       , fabric_tnd_hssl_atb_master_atdata_o28       =>  fabric_tnd_hssl_atb_master_atdata_o(27)
       , fabric_tnd_hssl_atb_master_atdata_o29       =>  fabric_tnd_hssl_atb_master_atdata_o(28)
       , fabric_tnd_hssl_atb_master_atdata_o30       =>  fabric_tnd_hssl_atb_master_atdata_o(29)
       , fabric_tnd_hssl_atb_master_atdata_o31       =>  fabric_tnd_hssl_atb_master_atdata_o(30)
       , fabric_tnd_hssl_atb_master_atdata_o32       =>  fabric_tnd_hssl_atb_master_atdata_o(31)
       , fabric_tnd_hssl_atb_master_atdata_o33       =>  fabric_tnd_hssl_atb_master_atdata_o(32)
       , fabric_tnd_hssl_atb_master_atdata_o34       =>  fabric_tnd_hssl_atb_master_atdata_o(33)
       , fabric_tnd_hssl_atb_master_atdata_o35       =>  fabric_tnd_hssl_atb_master_atdata_o(34)
       , fabric_tnd_hssl_atb_master_atdata_o36       =>  fabric_tnd_hssl_atb_master_atdata_o(35)
       , fabric_tnd_hssl_atb_master_atdata_o37       =>  fabric_tnd_hssl_atb_master_atdata_o(36)
       , fabric_tnd_hssl_atb_master_atdata_o38       =>  fabric_tnd_hssl_atb_master_atdata_o(37)
       , fabric_tnd_hssl_atb_master_atdata_o39       =>  fabric_tnd_hssl_atb_master_atdata_o(38)
       , fabric_tnd_hssl_atb_master_atdata_o40       =>  fabric_tnd_hssl_atb_master_atdata_o(39)
       , fabric_tnd_hssl_atb_master_atdata_o41       =>  fabric_tnd_hssl_atb_master_atdata_o(40)
       , fabric_tnd_hssl_atb_master_atdata_o42       =>  fabric_tnd_hssl_atb_master_atdata_o(41)
       , fabric_tnd_hssl_atb_master_atdata_o43       =>  fabric_tnd_hssl_atb_master_atdata_o(42)
       , fabric_tnd_hssl_atb_master_atdata_o44       =>  fabric_tnd_hssl_atb_master_atdata_o(43)
       , fabric_tnd_hssl_atb_master_atdata_o45       =>  fabric_tnd_hssl_atb_master_atdata_o(44)
       , fabric_tnd_hssl_atb_master_atdata_o46       =>  fabric_tnd_hssl_atb_master_atdata_o(45)
       , fabric_tnd_hssl_atb_master_atdata_o47       =>  fabric_tnd_hssl_atb_master_atdata_o(46)
       , fabric_tnd_hssl_atb_master_atdata_o48       =>  fabric_tnd_hssl_atb_master_atdata_o(47)
       , fabric_tnd_hssl_atb_master_atdata_o49       =>  fabric_tnd_hssl_atb_master_atdata_o(48)
       , fabric_tnd_hssl_atb_master_atdata_o50       =>  fabric_tnd_hssl_atb_master_atdata_o(49)
       , fabric_tnd_hssl_atb_master_atdata_o51       =>  fabric_tnd_hssl_atb_master_atdata_o(50)
       , fabric_tnd_hssl_atb_master_atdata_o52       =>  fabric_tnd_hssl_atb_master_atdata_o(51)
       , fabric_tnd_hssl_atb_master_atdata_o53       =>  fabric_tnd_hssl_atb_master_atdata_o(52)
       , fabric_tnd_hssl_atb_master_atdata_o54       =>  fabric_tnd_hssl_atb_master_atdata_o(53)
       , fabric_tnd_hssl_atb_master_atdata_o55       =>  fabric_tnd_hssl_atb_master_atdata_o(54)
       , fabric_tnd_hssl_atb_master_atdata_o56       =>  fabric_tnd_hssl_atb_master_atdata_o(55)
       , fabric_tnd_hssl_atb_master_atdata_o57       =>  fabric_tnd_hssl_atb_master_atdata_o(56)
       , fabric_tnd_hssl_atb_master_atdata_o58       =>  fabric_tnd_hssl_atb_master_atdata_o(57)
       , fabric_tnd_hssl_atb_master_atdata_o59       =>  fabric_tnd_hssl_atb_master_atdata_o(58)
       , fabric_tnd_hssl_atb_master_atdata_o60       =>  fabric_tnd_hssl_atb_master_atdata_o(59)
       , fabric_tnd_hssl_atb_master_atdata_o61       =>  fabric_tnd_hssl_atb_master_atdata_o(60)
       , fabric_tnd_hssl_atb_master_atdata_o62       =>  fabric_tnd_hssl_atb_master_atdata_o(61)
       , fabric_tnd_hssl_atb_master_atdata_o63       =>  fabric_tnd_hssl_atb_master_atdata_o(62)
       , fabric_tnd_hssl_atb_master_atdata_o64       =>  fabric_tnd_hssl_atb_master_atdata_o(63)
       , fabric_tnd_hssl_atb_master_atdata_o65       =>  fabric_tnd_hssl_atb_master_atdata_o(64)
       , fabric_tnd_hssl_atb_master_atdata_o66       =>  fabric_tnd_hssl_atb_master_atdata_o(65)
       , fabric_tnd_hssl_atb_master_atdata_o67       =>  fabric_tnd_hssl_atb_master_atdata_o(66)
       , fabric_tnd_hssl_atb_master_atdata_o68       =>  fabric_tnd_hssl_atb_master_atdata_o(67)
       , fabric_tnd_hssl_atb_master_atdata_o69       =>  fabric_tnd_hssl_atb_master_atdata_o(68)
       , fabric_tnd_hssl_atb_master_atdata_o70       =>  fabric_tnd_hssl_atb_master_atdata_o(69)
       , fabric_tnd_hssl_atb_master_atdata_o71       =>  fabric_tnd_hssl_atb_master_atdata_o(70)
       , fabric_tnd_hssl_atb_master_atdata_o72       =>  fabric_tnd_hssl_atb_master_atdata_o(71)
       , fabric_tnd_hssl_atb_master_atdata_o73       =>  fabric_tnd_hssl_atb_master_atdata_o(72)
       , fabric_tnd_hssl_atb_master_atdata_o74       =>  fabric_tnd_hssl_atb_master_atdata_o(73)
       , fabric_tnd_hssl_atb_master_atdata_o75       =>  fabric_tnd_hssl_atb_master_atdata_o(74)
       , fabric_tnd_hssl_atb_master_atdata_o76       =>  fabric_tnd_hssl_atb_master_atdata_o(75)
       , fabric_tnd_hssl_atb_master_atdata_o77       =>  fabric_tnd_hssl_atb_master_atdata_o(76)
       , fabric_tnd_hssl_atb_master_atdata_o78       =>  fabric_tnd_hssl_atb_master_atdata_o(77)
       , fabric_tnd_hssl_atb_master_atdata_o79       =>  fabric_tnd_hssl_atb_master_atdata_o(78)
       , fabric_tnd_hssl_atb_master_atdata_o80       =>  fabric_tnd_hssl_atb_master_atdata_o(79)
       , fabric_tnd_hssl_atb_master_atdata_o81       =>  fabric_tnd_hssl_atb_master_atdata_o(80)
       , fabric_tnd_hssl_atb_master_atdata_o82       =>  fabric_tnd_hssl_atb_master_atdata_o(81)
       , fabric_tnd_hssl_atb_master_atdata_o83       =>  fabric_tnd_hssl_atb_master_atdata_o(82)
       , fabric_tnd_hssl_atb_master_atdata_o84       =>  fabric_tnd_hssl_atb_master_atdata_o(83)
       , fabric_tnd_hssl_atb_master_atdata_o85       =>  fabric_tnd_hssl_atb_master_atdata_o(84)
       , fabric_tnd_hssl_atb_master_atdata_o86       =>  fabric_tnd_hssl_atb_master_atdata_o(85)
       , fabric_tnd_hssl_atb_master_atdata_o87       =>  fabric_tnd_hssl_atb_master_atdata_o(86)
       , fabric_tnd_hssl_atb_master_atdata_o88       =>  fabric_tnd_hssl_atb_master_atdata_o(87)
       , fabric_tnd_hssl_atb_master_atdata_o89       =>  fabric_tnd_hssl_atb_master_atdata_o(88)
       , fabric_tnd_hssl_atb_master_atdata_o90       =>  fabric_tnd_hssl_atb_master_atdata_o(89)
       , fabric_tnd_hssl_atb_master_atdata_o91       =>  fabric_tnd_hssl_atb_master_atdata_o(90)
       , fabric_tnd_hssl_atb_master_atdata_o92       =>  fabric_tnd_hssl_atb_master_atdata_o(91)
       , fabric_tnd_hssl_atb_master_atdata_o93       =>  fabric_tnd_hssl_atb_master_atdata_o(92)
       , fabric_tnd_hssl_atb_master_atdata_o94       =>  fabric_tnd_hssl_atb_master_atdata_o(93)
       , fabric_tnd_hssl_atb_master_atdata_o95       =>  fabric_tnd_hssl_atb_master_atdata_o(94)
       , fabric_tnd_hssl_atb_master_atdata_o96       =>  fabric_tnd_hssl_atb_master_atdata_o(95)
       , fabric_tnd_hssl_atb_master_atdata_o97       =>  fabric_tnd_hssl_atb_master_atdata_o(96)
       , fabric_tnd_hssl_atb_master_atdata_o98       =>  fabric_tnd_hssl_atb_master_atdata_o(97)
       , fabric_tnd_hssl_atb_master_atdata_o99       =>  fabric_tnd_hssl_atb_master_atdata_o(98)
       , fabric_tnd_hssl_atb_master_atdata_o100      =>  fabric_tnd_hssl_atb_master_atdata_o(99)
       , fabric_tnd_hssl_atb_master_atdata_o101      =>  fabric_tnd_hssl_atb_master_atdata_o(100)
       , fabric_tnd_hssl_atb_master_atdata_o102      =>  fabric_tnd_hssl_atb_master_atdata_o(101)
       , fabric_tnd_hssl_atb_master_atdata_o103      =>  fabric_tnd_hssl_atb_master_atdata_o(102)
       , fabric_tnd_hssl_atb_master_atdata_o104      =>  fabric_tnd_hssl_atb_master_atdata_o(103)
       , fabric_tnd_hssl_atb_master_atdata_o105      =>  fabric_tnd_hssl_atb_master_atdata_o(104)
       , fabric_tnd_hssl_atb_master_atdata_o106      =>  fabric_tnd_hssl_atb_master_atdata_o(105)
       , fabric_tnd_hssl_atb_master_atdata_o107      =>  fabric_tnd_hssl_atb_master_atdata_o(106)
       , fabric_tnd_hssl_atb_master_atdata_o108      =>  fabric_tnd_hssl_atb_master_atdata_o(107)
       , fabric_tnd_hssl_atb_master_atdata_o109      =>  fabric_tnd_hssl_atb_master_atdata_o(108)
       , fabric_tnd_hssl_atb_master_atdata_o110      =>  fabric_tnd_hssl_atb_master_atdata_o(109)
       , fabric_tnd_hssl_atb_master_atdata_o111      =>  fabric_tnd_hssl_atb_master_atdata_o(110)
       , fabric_tnd_hssl_atb_master_atdata_o112      =>  fabric_tnd_hssl_atb_master_atdata_o(111)
       , fabric_tnd_hssl_atb_master_atdata_o113      =>  fabric_tnd_hssl_atb_master_atdata_o(112)
       , fabric_tnd_hssl_atb_master_atdata_o114      =>  fabric_tnd_hssl_atb_master_atdata_o(113)
       , fabric_tnd_hssl_atb_master_atdata_o115      =>  fabric_tnd_hssl_atb_master_atdata_o(114)
       , fabric_tnd_hssl_atb_master_atdata_o116      =>  fabric_tnd_hssl_atb_master_atdata_o(115)
       , fabric_tnd_hssl_atb_master_atdata_o117      =>  fabric_tnd_hssl_atb_master_atdata_o(116)
       , fabric_tnd_hssl_atb_master_atdata_o118      =>  fabric_tnd_hssl_atb_master_atdata_o(117)
       , fabric_tnd_hssl_atb_master_atdata_o119      =>  fabric_tnd_hssl_atb_master_atdata_o(118)
       , fabric_tnd_hssl_atb_master_atdata_o120      =>  fabric_tnd_hssl_atb_master_atdata_o(119)
       , fabric_tnd_hssl_atb_master_atdata_o121      =>  fabric_tnd_hssl_atb_master_atdata_o(120)
       , fabric_tnd_hssl_atb_master_atdata_o122      =>  fabric_tnd_hssl_atb_master_atdata_o(121)
       , fabric_tnd_hssl_atb_master_atdata_o123      =>  fabric_tnd_hssl_atb_master_atdata_o(122)
       , fabric_tnd_hssl_atb_master_atdata_o124      =>  fabric_tnd_hssl_atb_master_atdata_o(123)
       , fabric_tnd_hssl_atb_master_atdata_o125      =>  fabric_tnd_hssl_atb_master_atdata_o(124)
       , fabric_tnd_hssl_atb_master_atdata_o126      =>  fabric_tnd_hssl_atb_master_atdata_o(125)
       , fabric_tnd_hssl_atb_master_atdata_o127      =>  fabric_tnd_hssl_atb_master_atdata_o(126)
       , fabric_tnd_hssl_atb_master_atdata_o128      =>  fabric_tnd_hssl_atb_master_atdata_o(127)
       , fabric_tnd_hssl_atb_master_atid_o1          =>  fabric_tnd_hssl_atb_master_atid_o(0)
       , fabric_tnd_hssl_atb_master_atid_o2          =>  fabric_tnd_hssl_atb_master_atid_o(1)
       , fabric_tnd_hssl_atb_master_atid_o3          =>  fabric_tnd_hssl_atb_master_atid_o(2)
       , fabric_tnd_hssl_atb_master_atid_o4          =>  fabric_tnd_hssl_atb_master_atid_o(3)
       , fabric_tnd_hssl_atb_master_atid_o5          =>  fabric_tnd_hssl_atb_master_atid_o(4)
       , fabric_tnd_hssl_atb_master_atid_o6          =>  fabric_tnd_hssl_atb_master_atid_o(5)
       , fabric_tnd_hssl_atb_master_atid_o7          =>  fabric_tnd_hssl_atb_master_atid_o(6)
       , fabric_tnd_hssl_atb_master_atvalid_o        =>  fabric_tnd_hssl_atb_master_atvalid_o
       , fabric_tnd_trace_clk_traceoutportintf_o     =>  fabric_tnd_trace_clk_traceoutportintf_o
       , fabric_tnd_trace_ctl_traceoutportintf_o     =>  fabric_tnd_trace_ctl_traceoutportintf_o
       , fabric_tnd_trace_data_traceoutportintf_o1   =>  fabric_tnd_trace_data_traceoutportintf_o(0)
       , fabric_tnd_trace_data_traceoutportintf_o2   =>  fabric_tnd_trace_data_traceoutportintf_o(1)
       , fabric_tnd_trace_data_traceoutportintf_o3   =>  fabric_tnd_trace_data_traceoutportintf_o(2)
       , fabric_tnd_trace_data_traceoutportintf_o4   =>  fabric_tnd_trace_data_traceoutportintf_o(3)
       , fabric_tnd_trace_data_traceoutportintf_o5   =>  fabric_tnd_trace_data_traceoutportintf_o(4)
       , fabric_tnd_trace_data_traceoutportintf_o6   =>  fabric_tnd_trace_data_traceoutportintf_o(5)
       , fabric_tnd_trace_data_traceoutportintf_o7   =>  fabric_tnd_trace_data_traceoutportintf_o(6)
       , fabric_tnd_trace_data_traceoutportintf_o8   =>  fabric_tnd_trace_data_traceoutportintf_o(7)
       , fabric_tnd_trace_data_traceoutportintf_o9   =>  fabric_tnd_trace_data_traceoutportintf_o(8)
       , fabric_tnd_trace_data_traceoutportintf_o10  =>  fabric_tnd_trace_data_traceoutportintf_o(9)
       , fabric_tnd_trace_data_traceoutportintf_o11  =>  fabric_tnd_trace_data_traceoutportintf_o(10)
       , fabric_tnd_trace_data_traceoutportintf_o12  =>  fabric_tnd_trace_data_traceoutportintf_o(11)
       , fabric_tnd_trace_data_traceoutportintf_o13  =>  fabric_tnd_trace_data_traceoutportintf_o(12)
       , fabric_tnd_trace_data_traceoutportintf_o14  =>  fabric_tnd_trace_data_traceoutportintf_o(13)
       , fabric_tnd_trace_data_traceoutportintf_o15  =>  fabric_tnd_trace_data_traceoutportintf_o(14)
       , fabric_tnd_trace_data_traceoutportintf_o16  =>  fabric_tnd_trace_data_traceoutportintf_o(15)
       , fabric_tnd_trace_data_traceoutportintf_o17  =>  fabric_tnd_trace_data_traceoutportintf_o(16)
       , fabric_tnd_trace_data_traceoutportintf_o18  =>  fabric_tnd_trace_data_traceoutportintf_o(17)
       , fabric_tnd_trace_data_traceoutportintf_o19  =>  fabric_tnd_trace_data_traceoutportintf_o(18)
       , fabric_tnd_trace_data_traceoutportintf_o20  =>  fabric_tnd_trace_data_traceoutportintf_o(19)
       , fabric_tnd_trace_data_traceoutportintf_o21  =>  fabric_tnd_trace_data_traceoutportintf_o(20)
       , fabric_tnd_trace_data_traceoutportintf_o22  =>  fabric_tnd_trace_data_traceoutportintf_o(21)
       , fabric_tnd_trace_data_traceoutportintf_o23  =>  fabric_tnd_trace_data_traceoutportintf_o(22)
       , fabric_tnd_trace_data_traceoutportintf_o24  =>  fabric_tnd_trace_data_traceoutportintf_o(23)
       , fabric_tnd_trace_data_traceoutportintf_o25  =>  fabric_tnd_trace_data_traceoutportintf_o(24)
       , fabric_tnd_trace_data_traceoutportintf_o26  =>  fabric_tnd_trace_data_traceoutportintf_o(25)
       , fabric_tnd_trace_data_traceoutportintf_o27  =>  fabric_tnd_trace_data_traceoutportintf_o(26)
       , fabric_tnd_trace_data_traceoutportintf_o28  =>  fabric_tnd_trace_data_traceoutportintf_o(27)
       , fabric_tnd_trace_data_traceoutportintf_o29  =>  fabric_tnd_trace_data_traceoutportintf_o(28)
       , fabric_tnd_trace_data_traceoutportintf_o30  =>  fabric_tnd_trace_data_traceoutportintf_o(29)
       , fabric_tnd_trace_data_traceoutportintf_o31  =>  fabric_tnd_trace_data_traceoutportintf_o(30)
       , fabric_tnd_trace_data_traceoutportintf_o32  =>  fabric_tnd_trace_data_traceoutportintf_o(31)
       , fabric_tsvalue_tsgen_fpga_o1                =>  fabric_tsvalue_tsgen_fpga_o(0)
       , fabric_tsvalue_tsgen_fpga_o2                =>  fabric_tsvalue_tsgen_fpga_o(1)
       , fabric_tsvalue_tsgen_fpga_o3                =>  fabric_tsvalue_tsgen_fpga_o(2)
       , fabric_tsvalue_tsgen_fpga_o4                =>  fabric_tsvalue_tsgen_fpga_o(3)
       , fabric_tsvalue_tsgen_fpga_o5                =>  fabric_tsvalue_tsgen_fpga_o(4)
       , fabric_tsvalue_tsgen_fpga_o6                =>  fabric_tsvalue_tsgen_fpga_o(5)
       , fabric_tsvalue_tsgen_fpga_o7                =>  fabric_tsvalue_tsgen_fpga_o(6)
       , fabric_tsvalue_tsgen_fpga_o8                =>  fabric_tsvalue_tsgen_fpga_o(7)
       , fabric_tsvalue_tsgen_fpga_o9                =>  fabric_tsvalue_tsgen_fpga_o(8)
       , fabric_tsvalue_tsgen_fpga_o10               =>  fabric_tsvalue_tsgen_fpga_o(9)
       , fabric_tsvalue_tsgen_fpga_o11               =>  fabric_tsvalue_tsgen_fpga_o(10)
       , fabric_tsvalue_tsgen_fpga_o12               =>  fabric_tsvalue_tsgen_fpga_o(11)
       , fabric_tsvalue_tsgen_fpga_o13               =>  fabric_tsvalue_tsgen_fpga_o(12)
       , fabric_tsvalue_tsgen_fpga_o14               =>  fabric_tsvalue_tsgen_fpga_o(13)
       , fabric_tsvalue_tsgen_fpga_o15               =>  fabric_tsvalue_tsgen_fpga_o(14)
       , fabric_tsvalue_tsgen_fpga_o16               =>  fabric_tsvalue_tsgen_fpga_o(15)
       , fabric_tsvalue_tsgen_fpga_o17               =>  fabric_tsvalue_tsgen_fpga_o(16)
       , fabric_tsvalue_tsgen_fpga_o18               =>  fabric_tsvalue_tsgen_fpga_o(17)
       , fabric_tsvalue_tsgen_fpga_o19               =>  fabric_tsvalue_tsgen_fpga_o(18)
       , fabric_tsvalue_tsgen_fpga_o20               =>  fabric_tsvalue_tsgen_fpga_o(19)
       , fabric_tsvalue_tsgen_fpga_o21               =>  fabric_tsvalue_tsgen_fpga_o(20)
       , fabric_tsvalue_tsgen_fpga_o22               =>  fabric_tsvalue_tsgen_fpga_o(21)
       , fabric_tsvalue_tsgen_fpga_o23               =>  fabric_tsvalue_tsgen_fpga_o(22)
       , fabric_tsvalue_tsgen_fpga_o24               =>  fabric_tsvalue_tsgen_fpga_o(23)
       , fabric_tsvalue_tsgen_fpga_o25               =>  fabric_tsvalue_tsgen_fpga_o(24)
       , fabric_tsvalue_tsgen_fpga_o26               =>  fabric_tsvalue_tsgen_fpga_o(25)
       , fabric_tsvalue_tsgen_fpga_o27               =>  fabric_tsvalue_tsgen_fpga_o(26)
       , fabric_tsvalue_tsgen_fpga_o28               =>  fabric_tsvalue_tsgen_fpga_o(27)
       , fabric_tsvalue_tsgen_fpga_o29               =>  fabric_tsvalue_tsgen_fpga_o(28)
       , fabric_tsvalue_tsgen_fpga_o30               =>  fabric_tsvalue_tsgen_fpga_o(29)
       , fabric_tsvalue_tsgen_fpga_o31               =>  fabric_tsvalue_tsgen_fpga_o(30)
       , fabric_tsvalue_tsgen_fpga_o32               =>  fabric_tsvalue_tsgen_fpga_o(31)
       , fabric_tsvalue_tsgen_fpga_o33               =>  fabric_tsvalue_tsgen_fpga_o(32)
       , fabric_tsvalue_tsgen_fpga_o34               =>  fabric_tsvalue_tsgen_fpga_o(33)
       , fabric_tsvalue_tsgen_fpga_o35               =>  fabric_tsvalue_tsgen_fpga_o(34)
       , fabric_tsvalue_tsgen_fpga_o36               =>  fabric_tsvalue_tsgen_fpga_o(35)
       , fabric_tsvalue_tsgen_fpga_o37               =>  fabric_tsvalue_tsgen_fpga_o(36)
       , fabric_tsvalue_tsgen_fpga_o38               =>  fabric_tsvalue_tsgen_fpga_o(37)
       , fabric_tsvalue_tsgen_fpga_o39               =>  fabric_tsvalue_tsgen_fpga_o(38)
       , fabric_tsvalue_tsgen_fpga_o40               =>  fabric_tsvalue_tsgen_fpga_o(39)
       , fabric_tsvalue_tsgen_fpga_o41               =>  fabric_tsvalue_tsgen_fpga_o(40)
       , fabric_tsvalue_tsgen_fpga_o42               =>  fabric_tsvalue_tsgen_fpga_o(41)
       , fabric_tsvalue_tsgen_fpga_o43               =>  fabric_tsvalue_tsgen_fpga_o(42)
       , fabric_tsvalue_tsgen_fpga_o44               =>  fabric_tsvalue_tsgen_fpga_o(43)
       , fabric_tsvalue_tsgen_fpga_o45               =>  fabric_tsvalue_tsgen_fpga_o(44)
       , fabric_tsvalue_tsgen_fpga_o46               =>  fabric_tsvalue_tsgen_fpga_o(45)
       , fabric_tsvalue_tsgen_fpga_o47               =>  fabric_tsvalue_tsgen_fpga_o(46)
       , fabric_tsvalue_tsgen_fpga_o48               =>  fabric_tsvalue_tsgen_fpga_o(47)
       , fabric_tsvalue_tsgen_fpga_o49               =>  fabric_tsvalue_tsgen_fpga_o(48)
       , fabric_tsvalue_tsgen_fpga_o50               =>  fabric_tsvalue_tsgen_fpga_o(49)
       , fabric_tsvalue_tsgen_fpga_o51               =>  fabric_tsvalue_tsgen_fpga_o(50)
       , fabric_tsvalue_tsgen_fpga_o52               =>  fabric_tsvalue_tsgen_fpga_o(51)
       , fabric_tsvalue_tsgen_fpga_o53               =>  fabric_tsvalue_tsgen_fpga_o(52)
       , fabric_tsvalue_tsgen_fpga_o54               =>  fabric_tsvalue_tsgen_fpga_o(53)
       , fabric_tsvalue_tsgen_fpga_o55               =>  fabric_tsvalue_tsgen_fpga_o(54)
       , fabric_tsvalue_tsgen_fpga_o56               =>  fabric_tsvalue_tsgen_fpga_o(55)
       , fabric_tsvalue_tsgen_fpga_o57               =>  fabric_tsvalue_tsgen_fpga_o(56)
       , fabric_tsvalue_tsgen_fpga_o58               =>  fabric_tsvalue_tsgen_fpga_o(57)
       , fabric_tsvalue_tsgen_fpga_o59               =>  fabric_tsvalue_tsgen_fpga_o(58)
       , fabric_tsvalue_tsgen_fpga_o60               =>  fabric_tsvalue_tsgen_fpga_o(59)
       , fabric_tsvalue_tsgen_fpga_o61               =>  fabric_tsvalue_tsgen_fpga_o(60)
       , fabric_tsvalue_tsgen_fpga_o62               =>  fabric_tsvalue_tsgen_fpga_o(61)
       , fabric_tsvalue_tsgen_fpga_o63               =>  fabric_tsvalue_tsgen_fpga_o(62)
       , fabric_tsvalue_tsgen_fpga_o64               =>  fabric_tsvalue_tsgen_fpga_o(63)
       , fabric_tnd_fpga_apb_master_prdata_i1        =>  fabric_tnd_fpga_apb_master_prdata_i(0)
       , fabric_tnd_fpga_apb_master_prdata_i2        =>  fabric_tnd_fpga_apb_master_prdata_i(1)
       , fabric_tnd_fpga_apb_master_prdata_i3        =>  fabric_tnd_fpga_apb_master_prdata_i(2)
       , fabric_tnd_fpga_apb_master_prdata_i4        =>  fabric_tnd_fpga_apb_master_prdata_i(3)
       , fabric_tnd_fpga_apb_master_prdata_i5        =>  fabric_tnd_fpga_apb_master_prdata_i(4)
       , fabric_tnd_fpga_apb_master_prdata_i6        =>  fabric_tnd_fpga_apb_master_prdata_i(5)
       , fabric_tnd_fpga_apb_master_prdata_i7        =>  fabric_tnd_fpga_apb_master_prdata_i(6)
       , fabric_tnd_fpga_apb_master_prdata_i8        =>  fabric_tnd_fpga_apb_master_prdata_i(7)
       , fabric_tnd_fpga_apb_master_prdata_i9        =>  fabric_tnd_fpga_apb_master_prdata_i(8)
       , fabric_tnd_fpga_apb_master_prdata_i10       =>  fabric_tnd_fpga_apb_master_prdata_i(9)
       , fabric_tnd_fpga_apb_master_prdata_i11       =>  fabric_tnd_fpga_apb_master_prdata_i(10)
       , fabric_tnd_fpga_apb_master_prdata_i12       =>  fabric_tnd_fpga_apb_master_prdata_i(11)
       , fabric_tnd_fpga_apb_master_prdata_i13       =>  fabric_tnd_fpga_apb_master_prdata_i(12)
       , fabric_tnd_fpga_apb_master_prdata_i14       =>  fabric_tnd_fpga_apb_master_prdata_i(13)
       , fabric_tnd_fpga_apb_master_prdata_i15       =>  fabric_tnd_fpga_apb_master_prdata_i(14)
       , fabric_tnd_fpga_apb_master_prdata_i16       =>  fabric_tnd_fpga_apb_master_prdata_i(15)
       , fabric_tnd_fpga_apb_master_prdata_i17       =>  fabric_tnd_fpga_apb_master_prdata_i(16)
       , fabric_tnd_fpga_apb_master_prdata_i18       =>  fabric_tnd_fpga_apb_master_prdata_i(17)
       , fabric_tnd_fpga_apb_master_prdata_i19       =>  fabric_tnd_fpga_apb_master_prdata_i(18)
       , fabric_tnd_fpga_apb_master_prdata_i20       =>  fabric_tnd_fpga_apb_master_prdata_i(19)
       , fabric_tnd_fpga_apb_master_prdata_i21       =>  fabric_tnd_fpga_apb_master_prdata_i(20)
       , fabric_tnd_fpga_apb_master_prdata_i22       =>  fabric_tnd_fpga_apb_master_prdata_i(21)
       , fabric_tnd_fpga_apb_master_prdata_i23       =>  fabric_tnd_fpga_apb_master_prdata_i(22)
       , fabric_tnd_fpga_apb_master_prdata_i24       =>  fabric_tnd_fpga_apb_master_prdata_i(23)
       , fabric_tnd_fpga_apb_master_prdata_i25       =>  fabric_tnd_fpga_apb_master_prdata_i(24)
       , fabric_tnd_fpga_apb_master_prdata_i26       =>  fabric_tnd_fpga_apb_master_prdata_i(25)
       , fabric_tnd_fpga_apb_master_prdata_i27       =>  fabric_tnd_fpga_apb_master_prdata_i(26)
       , fabric_tnd_fpga_apb_master_prdata_i28       =>  fabric_tnd_fpga_apb_master_prdata_i(27)
       , fabric_tnd_fpga_apb_master_prdata_i29       =>  fabric_tnd_fpga_apb_master_prdata_i(28)
       , fabric_tnd_fpga_apb_master_prdata_i30       =>  fabric_tnd_fpga_apb_master_prdata_i(29)
       , fabric_tnd_fpga_apb_master_prdata_i31       =>  fabric_tnd_fpga_apb_master_prdata_i(30)
       , fabric_tnd_fpga_apb_master_prdata_i32       =>  fabric_tnd_fpga_apb_master_prdata_i(31)
       , fabric_tnd_fpga_apb_master_pready_i         =>  fabric_tnd_fpga_apb_master_pready_i
       , fabric_tnd_fpga_apb_master_pslverr_i        =>  fabric_tnd_fpga_apb_master_pslverr_i
       , fabric_tnd_fpga_atb_master_afready_i        =>  fabric_tnd_fpga_atb_master_afready_i
       , fabric_tnd_fpga_atb_master_atbytes_i1       =>  fabric_tnd_fpga_atb_master_atbytes_i(0)
       , fabric_tnd_fpga_atb_master_atbytes_i2       =>  fabric_tnd_fpga_atb_master_atbytes_i(1)
       , fabric_tnd_fpga_atb_master_atbytes_i3       =>  fabric_tnd_fpga_atb_master_atbytes_i(2)
       , fabric_tnd_fpga_atb_master_atbytes_i4       =>  fabric_tnd_fpga_atb_master_atbytes_i(3)
       , fabric_tnd_fpga_atb_master_atdata_i1        =>  fabric_tnd_fpga_atb_master_atdata_i(0)
       , fabric_tnd_fpga_atb_master_atdata_i2        =>  fabric_tnd_fpga_atb_master_atdata_i(1)
       , fabric_tnd_fpga_atb_master_atdata_i3        =>  fabric_tnd_fpga_atb_master_atdata_i(2)
       , fabric_tnd_fpga_atb_master_atdata_i4        =>  fabric_tnd_fpga_atb_master_atdata_i(3)
       , fabric_tnd_fpga_atb_master_atdata_i5        =>  fabric_tnd_fpga_atb_master_atdata_i(4)
       , fabric_tnd_fpga_atb_master_atdata_i6        =>  fabric_tnd_fpga_atb_master_atdata_i(5)
       , fabric_tnd_fpga_atb_master_atdata_i7        =>  fabric_tnd_fpga_atb_master_atdata_i(6)
       , fabric_tnd_fpga_atb_master_atdata_i8        =>  fabric_tnd_fpga_atb_master_atdata_i(7)
       , fabric_tnd_fpga_atb_master_atdata_i9        =>  fabric_tnd_fpga_atb_master_atdata_i(8)
       , fabric_tnd_fpga_atb_master_atdata_i10       =>  fabric_tnd_fpga_atb_master_atdata_i(9)
       , fabric_tnd_fpga_atb_master_atdata_i11       =>  fabric_tnd_fpga_atb_master_atdata_i(10)
       , fabric_tnd_fpga_atb_master_atdata_i12       =>  fabric_tnd_fpga_atb_master_atdata_i(11)
       , fabric_tnd_fpga_atb_master_atdata_i13       =>  fabric_tnd_fpga_atb_master_atdata_i(12)
       , fabric_tnd_fpga_atb_master_atdata_i14       =>  fabric_tnd_fpga_atb_master_atdata_i(13)
       , fabric_tnd_fpga_atb_master_atdata_i15       =>  fabric_tnd_fpga_atb_master_atdata_i(14)
       , fabric_tnd_fpga_atb_master_atdata_i16       =>  fabric_tnd_fpga_atb_master_atdata_i(15)
       , fabric_tnd_fpga_atb_master_atdata_i17       =>  fabric_tnd_fpga_atb_master_atdata_i(16)
       , fabric_tnd_fpga_atb_master_atdata_i18       =>  fabric_tnd_fpga_atb_master_atdata_i(17)
       , fabric_tnd_fpga_atb_master_atdata_i19       =>  fabric_tnd_fpga_atb_master_atdata_i(18)
       , fabric_tnd_fpga_atb_master_atdata_i20       =>  fabric_tnd_fpga_atb_master_atdata_i(19)
       , fabric_tnd_fpga_atb_master_atdata_i21       =>  fabric_tnd_fpga_atb_master_atdata_i(20)
       , fabric_tnd_fpga_atb_master_atdata_i22       =>  fabric_tnd_fpga_atb_master_atdata_i(21)
       , fabric_tnd_fpga_atb_master_atdata_i23       =>  fabric_tnd_fpga_atb_master_atdata_i(22)
       , fabric_tnd_fpga_atb_master_atdata_i24       =>  fabric_tnd_fpga_atb_master_atdata_i(23)
       , fabric_tnd_fpga_atb_master_atdata_i25       =>  fabric_tnd_fpga_atb_master_atdata_i(24)
       , fabric_tnd_fpga_atb_master_atdata_i26       =>  fabric_tnd_fpga_atb_master_atdata_i(25)
       , fabric_tnd_fpga_atb_master_atdata_i27       =>  fabric_tnd_fpga_atb_master_atdata_i(26)
       , fabric_tnd_fpga_atb_master_atdata_i28       =>  fabric_tnd_fpga_atb_master_atdata_i(27)
       , fabric_tnd_fpga_atb_master_atdata_i29       =>  fabric_tnd_fpga_atb_master_atdata_i(28)
       , fabric_tnd_fpga_atb_master_atdata_i30       =>  fabric_tnd_fpga_atb_master_atdata_i(29)
       , fabric_tnd_fpga_atb_master_atdata_i31       =>  fabric_tnd_fpga_atb_master_atdata_i(30)
       , fabric_tnd_fpga_atb_master_atdata_i32       =>  fabric_tnd_fpga_atb_master_atdata_i(31)
       , fabric_tnd_fpga_atb_master_atdata_i33       =>  fabric_tnd_fpga_atb_master_atdata_i(32)
       , fabric_tnd_fpga_atb_master_atdata_i34       =>  fabric_tnd_fpga_atb_master_atdata_i(33)
       , fabric_tnd_fpga_atb_master_atdata_i35       =>  fabric_tnd_fpga_atb_master_atdata_i(34)
       , fabric_tnd_fpga_atb_master_atdata_i36       =>  fabric_tnd_fpga_atb_master_atdata_i(35)
       , fabric_tnd_fpga_atb_master_atdata_i37       =>  fabric_tnd_fpga_atb_master_atdata_i(36)
       , fabric_tnd_fpga_atb_master_atdata_i38       =>  fabric_tnd_fpga_atb_master_atdata_i(37)
       , fabric_tnd_fpga_atb_master_atdata_i39       =>  fabric_tnd_fpga_atb_master_atdata_i(38)
       , fabric_tnd_fpga_atb_master_atdata_i40       =>  fabric_tnd_fpga_atb_master_atdata_i(39)
       , fabric_tnd_fpga_atb_master_atdata_i41       =>  fabric_tnd_fpga_atb_master_atdata_i(40)
       , fabric_tnd_fpga_atb_master_atdata_i42       =>  fabric_tnd_fpga_atb_master_atdata_i(41)
       , fabric_tnd_fpga_atb_master_atdata_i43       =>  fabric_tnd_fpga_atb_master_atdata_i(42)
       , fabric_tnd_fpga_atb_master_atdata_i44       =>  fabric_tnd_fpga_atb_master_atdata_i(43)
       , fabric_tnd_fpga_atb_master_atdata_i45       =>  fabric_tnd_fpga_atb_master_atdata_i(44)
       , fabric_tnd_fpga_atb_master_atdata_i46       =>  fabric_tnd_fpga_atb_master_atdata_i(45)
       , fabric_tnd_fpga_atb_master_atdata_i47       =>  fabric_tnd_fpga_atb_master_atdata_i(46)
       , fabric_tnd_fpga_atb_master_atdata_i48       =>  fabric_tnd_fpga_atb_master_atdata_i(47)
       , fabric_tnd_fpga_atb_master_atdata_i49       =>  fabric_tnd_fpga_atb_master_atdata_i(48)
       , fabric_tnd_fpga_atb_master_atdata_i50       =>  fabric_tnd_fpga_atb_master_atdata_i(49)
       , fabric_tnd_fpga_atb_master_atdata_i51       =>  fabric_tnd_fpga_atb_master_atdata_i(50)
       , fabric_tnd_fpga_atb_master_atdata_i52       =>  fabric_tnd_fpga_atb_master_atdata_i(51)
       , fabric_tnd_fpga_atb_master_atdata_i53       =>  fabric_tnd_fpga_atb_master_atdata_i(52)
       , fabric_tnd_fpga_atb_master_atdata_i54       =>  fabric_tnd_fpga_atb_master_atdata_i(53)
       , fabric_tnd_fpga_atb_master_atdata_i55       =>  fabric_tnd_fpga_atb_master_atdata_i(54)
       , fabric_tnd_fpga_atb_master_atdata_i56       =>  fabric_tnd_fpga_atb_master_atdata_i(55)
       , fabric_tnd_fpga_atb_master_atdata_i57       =>  fabric_tnd_fpga_atb_master_atdata_i(56)
       , fabric_tnd_fpga_atb_master_atdata_i58       =>  fabric_tnd_fpga_atb_master_atdata_i(57)
       , fabric_tnd_fpga_atb_master_atdata_i59       =>  fabric_tnd_fpga_atb_master_atdata_i(58)
       , fabric_tnd_fpga_atb_master_atdata_i60       =>  fabric_tnd_fpga_atb_master_atdata_i(59)
       , fabric_tnd_fpga_atb_master_atdata_i61       =>  fabric_tnd_fpga_atb_master_atdata_i(60)
       , fabric_tnd_fpga_atb_master_atdata_i62       =>  fabric_tnd_fpga_atb_master_atdata_i(61)
       , fabric_tnd_fpga_atb_master_atdata_i63       =>  fabric_tnd_fpga_atb_master_atdata_i(62)
       , fabric_tnd_fpga_atb_master_atdata_i64       =>  fabric_tnd_fpga_atb_master_atdata_i(63)
       , fabric_tnd_fpga_atb_master_atdata_i65       =>  fabric_tnd_fpga_atb_master_atdata_i(64)
       , fabric_tnd_fpga_atb_master_atdata_i66       =>  fabric_tnd_fpga_atb_master_atdata_i(65)
       , fabric_tnd_fpga_atb_master_atdata_i67       =>  fabric_tnd_fpga_atb_master_atdata_i(66)
       , fabric_tnd_fpga_atb_master_atdata_i68       =>  fabric_tnd_fpga_atb_master_atdata_i(67)
       , fabric_tnd_fpga_atb_master_atdata_i69       =>  fabric_tnd_fpga_atb_master_atdata_i(68)
       , fabric_tnd_fpga_atb_master_atdata_i70       =>  fabric_tnd_fpga_atb_master_atdata_i(69)
       , fabric_tnd_fpga_atb_master_atdata_i71       =>  fabric_tnd_fpga_atb_master_atdata_i(70)
       , fabric_tnd_fpga_atb_master_atdata_i72       =>  fabric_tnd_fpga_atb_master_atdata_i(71)
       , fabric_tnd_fpga_atb_master_atdata_i73       =>  fabric_tnd_fpga_atb_master_atdata_i(72)
       , fabric_tnd_fpga_atb_master_atdata_i74       =>  fabric_tnd_fpga_atb_master_atdata_i(73)
       , fabric_tnd_fpga_atb_master_atdata_i75       =>  fabric_tnd_fpga_atb_master_atdata_i(74)
       , fabric_tnd_fpga_atb_master_atdata_i76       =>  fabric_tnd_fpga_atb_master_atdata_i(75)
       , fabric_tnd_fpga_atb_master_atdata_i77       =>  fabric_tnd_fpga_atb_master_atdata_i(76)
       , fabric_tnd_fpga_atb_master_atdata_i78       =>  fabric_tnd_fpga_atb_master_atdata_i(77)
       , fabric_tnd_fpga_atb_master_atdata_i79       =>  fabric_tnd_fpga_atb_master_atdata_i(78)
       , fabric_tnd_fpga_atb_master_atdata_i80       =>  fabric_tnd_fpga_atb_master_atdata_i(79)
       , fabric_tnd_fpga_atb_master_atdata_i81       =>  fabric_tnd_fpga_atb_master_atdata_i(80)
       , fabric_tnd_fpga_atb_master_atdata_i82       =>  fabric_tnd_fpga_atb_master_atdata_i(81)
       , fabric_tnd_fpga_atb_master_atdata_i83       =>  fabric_tnd_fpga_atb_master_atdata_i(82)
       , fabric_tnd_fpga_atb_master_atdata_i84       =>  fabric_tnd_fpga_atb_master_atdata_i(83)
       , fabric_tnd_fpga_atb_master_atdata_i85       =>  fabric_tnd_fpga_atb_master_atdata_i(84)
       , fabric_tnd_fpga_atb_master_atdata_i86       =>  fabric_tnd_fpga_atb_master_atdata_i(85)
       , fabric_tnd_fpga_atb_master_atdata_i87       =>  fabric_tnd_fpga_atb_master_atdata_i(86)
       , fabric_tnd_fpga_atb_master_atdata_i88       =>  fabric_tnd_fpga_atb_master_atdata_i(87)
       , fabric_tnd_fpga_atb_master_atdata_i89       =>  fabric_tnd_fpga_atb_master_atdata_i(88)
       , fabric_tnd_fpga_atb_master_atdata_i90       =>  fabric_tnd_fpga_atb_master_atdata_i(89)
       , fabric_tnd_fpga_atb_master_atdata_i91       =>  fabric_tnd_fpga_atb_master_atdata_i(90)
       , fabric_tnd_fpga_atb_master_atdata_i92       =>  fabric_tnd_fpga_atb_master_atdata_i(91)
       , fabric_tnd_fpga_atb_master_atdata_i93       =>  fabric_tnd_fpga_atb_master_atdata_i(92)
       , fabric_tnd_fpga_atb_master_atdata_i94       =>  fabric_tnd_fpga_atb_master_atdata_i(93)
       , fabric_tnd_fpga_atb_master_atdata_i95       =>  fabric_tnd_fpga_atb_master_atdata_i(94)
       , fabric_tnd_fpga_atb_master_atdata_i96       =>  fabric_tnd_fpga_atb_master_atdata_i(95)
       , fabric_tnd_fpga_atb_master_atdata_i97       =>  fabric_tnd_fpga_atb_master_atdata_i(96)
       , fabric_tnd_fpga_atb_master_atdata_i98       =>  fabric_tnd_fpga_atb_master_atdata_i(97)
       , fabric_tnd_fpga_atb_master_atdata_i99       =>  fabric_tnd_fpga_atb_master_atdata_i(98)
       , fabric_tnd_fpga_atb_master_atdata_i100      =>  fabric_tnd_fpga_atb_master_atdata_i(99)
       , fabric_tnd_fpga_atb_master_atdata_i101      =>  fabric_tnd_fpga_atb_master_atdata_i(100)
       , fabric_tnd_fpga_atb_master_atdata_i102      =>  fabric_tnd_fpga_atb_master_atdata_i(101)
       , fabric_tnd_fpga_atb_master_atdata_i103      =>  fabric_tnd_fpga_atb_master_atdata_i(102)
       , fabric_tnd_fpga_atb_master_atdata_i104      =>  fabric_tnd_fpga_atb_master_atdata_i(103)
       , fabric_tnd_fpga_atb_master_atdata_i105      =>  fabric_tnd_fpga_atb_master_atdata_i(104)
       , fabric_tnd_fpga_atb_master_atdata_i106      =>  fabric_tnd_fpga_atb_master_atdata_i(105)
       , fabric_tnd_fpga_atb_master_atdata_i107      =>  fabric_tnd_fpga_atb_master_atdata_i(106)
       , fabric_tnd_fpga_atb_master_atdata_i108      =>  fabric_tnd_fpga_atb_master_atdata_i(107)
       , fabric_tnd_fpga_atb_master_atdata_i109      =>  fabric_tnd_fpga_atb_master_atdata_i(108)
       , fabric_tnd_fpga_atb_master_atdata_i110      =>  fabric_tnd_fpga_atb_master_atdata_i(109)
       , fabric_tnd_fpga_atb_master_atdata_i111      =>  fabric_tnd_fpga_atb_master_atdata_i(110)
       , fabric_tnd_fpga_atb_master_atdata_i112      =>  fabric_tnd_fpga_atb_master_atdata_i(111)
       , fabric_tnd_fpga_atb_master_atdata_i113      =>  fabric_tnd_fpga_atb_master_atdata_i(112)
       , fabric_tnd_fpga_atb_master_atdata_i114      =>  fabric_tnd_fpga_atb_master_atdata_i(113)
       , fabric_tnd_fpga_atb_master_atdata_i115      =>  fabric_tnd_fpga_atb_master_atdata_i(114)
       , fabric_tnd_fpga_atb_master_atdata_i116      =>  fabric_tnd_fpga_atb_master_atdata_i(115)
       , fabric_tnd_fpga_atb_master_atdata_i117      =>  fabric_tnd_fpga_atb_master_atdata_i(116)
       , fabric_tnd_fpga_atb_master_atdata_i118      =>  fabric_tnd_fpga_atb_master_atdata_i(117)
       , fabric_tnd_fpga_atb_master_atdata_i119      =>  fabric_tnd_fpga_atb_master_atdata_i(118)
       , fabric_tnd_fpga_atb_master_atdata_i120      =>  fabric_tnd_fpga_atb_master_atdata_i(119)
       , fabric_tnd_fpga_atb_master_atdata_i121      =>  fabric_tnd_fpga_atb_master_atdata_i(120)
       , fabric_tnd_fpga_atb_master_atdata_i122      =>  fabric_tnd_fpga_atb_master_atdata_i(121)
       , fabric_tnd_fpga_atb_master_atdata_i123      =>  fabric_tnd_fpga_atb_master_atdata_i(122)
       , fabric_tnd_fpga_atb_master_atdata_i124      =>  fabric_tnd_fpga_atb_master_atdata_i(123)
       , fabric_tnd_fpga_atb_master_atdata_i125      =>  fabric_tnd_fpga_atb_master_atdata_i(124)
       , fabric_tnd_fpga_atb_master_atdata_i126      =>  fabric_tnd_fpga_atb_master_atdata_i(125)
       , fabric_tnd_fpga_atb_master_atdata_i127      =>  fabric_tnd_fpga_atb_master_atdata_i(126)
       , fabric_tnd_fpga_atb_master_atdata_i128      =>  fabric_tnd_fpga_atb_master_atdata_i(127)
       , fabric_tnd_fpga_atb_master_atid_i1          =>  fabric_tnd_fpga_atb_master_atid_i(0)
       , fabric_tnd_fpga_atb_master_atid_i2          =>  fabric_tnd_fpga_atb_master_atid_i(1)
       , fabric_tnd_fpga_atb_master_atid_i3          =>  fabric_tnd_fpga_atb_master_atid_i(2)
       , fabric_tnd_fpga_atb_master_atid_i4          =>  fabric_tnd_fpga_atb_master_atid_i(3)
       , fabric_tnd_fpga_atb_master_atid_i5          =>  fabric_tnd_fpga_atb_master_atid_i(4)
       , fabric_tnd_fpga_atb_master_atid_i6          =>  fabric_tnd_fpga_atb_master_atid_i(5)
       , fabric_tnd_fpga_atb_master_atid_i7          =>  fabric_tnd_fpga_atb_master_atid_i(6)
       , fabric_tnd_fpga_atb_master_atvalid_i        =>  fabric_tnd_fpga_atb_master_atvalid_i
       , fabric_tnd_hssl_apb_master_prdata_i1        =>  fabric_tnd_hssl_apb_master_prdata_i(0)
       , fabric_tnd_hssl_apb_master_prdata_i2        =>  fabric_tnd_hssl_apb_master_prdata_i(1)
       , fabric_tnd_hssl_apb_master_prdata_i3        =>  fabric_tnd_hssl_apb_master_prdata_i(2)
       , fabric_tnd_hssl_apb_master_prdata_i4        =>  fabric_tnd_hssl_apb_master_prdata_i(3)
       , fabric_tnd_hssl_apb_master_prdata_i5        =>  fabric_tnd_hssl_apb_master_prdata_i(4)
       , fabric_tnd_hssl_apb_master_prdata_i6        =>  fabric_tnd_hssl_apb_master_prdata_i(5)
       , fabric_tnd_hssl_apb_master_prdata_i7        =>  fabric_tnd_hssl_apb_master_prdata_i(6)
       , fabric_tnd_hssl_apb_master_prdata_i8        =>  fabric_tnd_hssl_apb_master_prdata_i(7)
       , fabric_tnd_hssl_apb_master_prdata_i9        =>  fabric_tnd_hssl_apb_master_prdata_i(8)
       , fabric_tnd_hssl_apb_master_prdata_i10       =>  fabric_tnd_hssl_apb_master_prdata_i(9)
       , fabric_tnd_hssl_apb_master_prdata_i11       =>  fabric_tnd_hssl_apb_master_prdata_i(10)
       , fabric_tnd_hssl_apb_master_prdata_i12       =>  fabric_tnd_hssl_apb_master_prdata_i(11)
       , fabric_tnd_hssl_apb_master_prdata_i13       =>  fabric_tnd_hssl_apb_master_prdata_i(12)
       , fabric_tnd_hssl_apb_master_prdata_i14       =>  fabric_tnd_hssl_apb_master_prdata_i(13)
       , fabric_tnd_hssl_apb_master_prdata_i15       =>  fabric_tnd_hssl_apb_master_prdata_i(14)
       , fabric_tnd_hssl_apb_master_prdata_i16       =>  fabric_tnd_hssl_apb_master_prdata_i(15)
       , fabric_tnd_hssl_apb_master_prdata_i17       =>  fabric_tnd_hssl_apb_master_prdata_i(16)
       , fabric_tnd_hssl_apb_master_prdata_i18       =>  fabric_tnd_hssl_apb_master_prdata_i(17)
       , fabric_tnd_hssl_apb_master_prdata_i19       =>  fabric_tnd_hssl_apb_master_prdata_i(18)
       , fabric_tnd_hssl_apb_master_prdata_i20       =>  fabric_tnd_hssl_apb_master_prdata_i(19)
       , fabric_tnd_hssl_apb_master_prdata_i21       =>  fabric_tnd_hssl_apb_master_prdata_i(20)
       , fabric_tnd_hssl_apb_master_prdata_i22       =>  fabric_tnd_hssl_apb_master_prdata_i(21)
       , fabric_tnd_hssl_apb_master_prdata_i23       =>  fabric_tnd_hssl_apb_master_prdata_i(22)
       , fabric_tnd_hssl_apb_master_prdata_i24       =>  fabric_tnd_hssl_apb_master_prdata_i(23)
       , fabric_tnd_hssl_apb_master_prdata_i25       =>  fabric_tnd_hssl_apb_master_prdata_i(24)
       , fabric_tnd_hssl_apb_master_prdata_i26       =>  fabric_tnd_hssl_apb_master_prdata_i(25)
       , fabric_tnd_hssl_apb_master_prdata_i27       =>  fabric_tnd_hssl_apb_master_prdata_i(26)
       , fabric_tnd_hssl_apb_master_prdata_i28       =>  fabric_tnd_hssl_apb_master_prdata_i(27)
       , fabric_tnd_hssl_apb_master_prdata_i29       =>  fabric_tnd_hssl_apb_master_prdata_i(28)
       , fabric_tnd_hssl_apb_master_prdata_i30       =>  fabric_tnd_hssl_apb_master_prdata_i(29)
       , fabric_tnd_hssl_apb_master_prdata_i31       =>  fabric_tnd_hssl_apb_master_prdata_i(30)
       , fabric_tnd_hssl_apb_master_prdata_i32       =>  fabric_tnd_hssl_apb_master_prdata_i(31)
       , fabric_tnd_hssl_apb_master_pready_i         =>  fabric_tnd_hssl_apb_master_pready_i
       , fabric_tnd_hssl_apb_master_pslverr_i        =>  fabric_tnd_hssl_apb_master_pslverr_i
       , fabric_tnd_hssl_atb_master_afvalid_i        =>  fabric_tnd_hssl_atb_master_afvalid_i
       , fabric_tnd_hssl_atb_master_atready_i        =>  fabric_tnd_hssl_atb_master_atready_i
       , fabric_tnd_hssl_atb_master_syncreq_i        =>  fabric_tnd_hssl_atb_master_syncreq_i
       , fabric_watchdog0_signal_0_o                 =>  fabric_watchdog0_signal_0_o
       , fabric_watchdog0_signal_1_o                 =>  fabric_watchdog0_signal_1_o
       , fabric_watchdog1_signal_0_o                 =>  fabric_watchdog1_signal_0_o
       , fabric_watchdog1_signal_1_o                 =>  fabric_watchdog1_signal_1_o
       , fabric_watchdog2_signal_0_o                 =>  fabric_watchdog2_signal_0_o
       , fabric_watchdog2_signal_1_o                 =>  fabric_watchdog2_signal_1_o
       , fabric_watchdog3_signal_0_o                 =>  fabric_watchdog3_signal_0_o
       , fabric_watchdog3_signal_1_o                 =>  fabric_watchdog3_signal_1_o
       , fabric_tst_pll_lock_o1                      =>  fabric_tst_pll_lock_o(0)
       , fabric_tst_pll_lock_o2                      =>  fabric_tst_pll_lock_o(1)
       , fabric_tst_pll_lock_o3                      =>  fabric_tst_pll_lock_o(2)
       , fabric_tst_pll_lock_o4                      =>  fabric_tst_pll_lock_o(3)
       , fabric_tst_pll_lock_o5                      =>  fabric_tst_pll_lock_o(4)
       , fabric_tst_pll_lock_o6                      =>  fabric_tst_pll_lock_o(5)
       , fabric_tst_pll_lock_o7                      =>  fabric_tst_pll_lock_o(6)
       , fabric_soc_mon_sensor_alarm_o               =>  fabric_soc_mon_sensor_alarm_o
       , fabric_erom_fpga_cpu0_dbgen_i               =>  fabric_erom_fpga_cpu0_dbgen_i
       , fabric_erom_fpga_cpu0_hiden_i               =>  fabric_erom_fpga_cpu0_hiden_i
       , fabric_erom_fpga_cpu0_hniden_i              =>  fabric_erom_fpga_cpu0_hniden_i
       , fabric_erom_fpga_cpu0_niden_i               =>  fabric_erom_fpga_cpu0_niden_i
       , fabric_erom_fpga_cpu1_dbgen_i               =>  fabric_erom_fpga_cpu1_dbgen_i
       , fabric_erom_fpga_cpu1_hiden_i               =>  fabric_erom_fpga_cpu1_hiden_i
       , fabric_erom_fpga_cpu1_hniden_i              =>  fabric_erom_fpga_cpu1_hniden_i
       , fabric_erom_fpga_cpu1_niden_i               =>  fabric_erom_fpga_cpu1_niden_i
       , fabric_erom_fpga_cpu2_dbgen_i               =>  fabric_erom_fpga_cpu2_dbgen_i
       , fabric_erom_fpga_cpu2_hiden_i               =>  fabric_erom_fpga_cpu2_hiden_i
       , fabric_erom_fpga_cpu2_hniden_i              =>  fabric_erom_fpga_cpu2_hniden_i
       , fabric_erom_fpga_cpu2_niden_i               =>  fabric_erom_fpga_cpu2_niden_i
       , fabric_erom_fpga_cpu3_dbgen_i               =>  fabric_erom_fpga_cpu3_dbgen_i
       , fabric_erom_fpga_cpu3_hiden_i               =>  fabric_erom_fpga_cpu3_hiden_i
       , fabric_erom_fpga_cpu3_hniden_i              =>  fabric_erom_fpga_cpu3_hniden_i
       , fabric_erom_fpga_cpu3_niden_i               =>  fabric_erom_fpga_cpu3_niden_i
       , fabric_erom_fpga_cs_dbgen_i                 =>  fabric_erom_fpga_cs_dbgen_i
       , fabric_erom_fpga_cs_niden_i                 =>  fabric_erom_fpga_cs_niden_i
       , fabric_erom_fpga_cs_deviceen_i              =>  fabric_erom_fpga_cs_deviceen_i
       , fabric_erom_fpga_cs_rst_n_i                 =>  fabric_erom_fpga_cs_rst_n_i
       , fabric_erom_fpga_debug_en_i                 =>  fabric_erom_fpga_debug_en_i
       , fabric_enable_TMR_i1                        =>  fabric_enable_TMR_i(0)
       , fabric_enable_TMR_i2                        =>  fabric_enable_TMR_i(1)
       , fabric_enable_TMR_i3                        =>  fabric_enable_TMR_i(2)
);
end NX_RTL;

-- =================================================================================================
--   NX_BD definition                                                                   2018/06/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_BD is
generic (
    mode : string := "local_lowskew"
);
port (
    I : in  std_logic;
    O : out std_logic
);
end NX_BD;

-- =================================================================================================
--   NX_CY definition                                                                   2017/09/19
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_CY is
generic (
    add_carry  : integer := 0      -- 0: low - 1: high - 2: propagate
);
port (
    A1 : in  std_logic;
    A2 : in  std_logic;
    A3 : in  std_logic;
    A4 : in  std_logic;
    B1 : in  std_logic;
    B2 : in  std_logic;
    B3 : in  std_logic;
    B4 : in  std_logic;
    CI : in  std_logic;
    CO : out std_logic;
    S1 : out std_logic;
    S2 : out std_logic;
    S3 : out std_logic;
    S4 : out std_logic
);
end NX_CY;

-- =================================================================================================
--   NX_ECC definition                                                                  2020/05/12
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_ECC is
    port(
	CKD : in std_logic;
	CHK : in std_logic;
	COR : out std_logic;
	ERR : out std_logic
    );
end NX_ECC;
-- =================================================================================================
--   NX_LUT definition                                                                  2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_LUT is
generic (
    lut_table : bit_vector(15 downto 0) := B"0000000000000000" -- truthTable t15 ... t0
);
port (
    I1 : in  std_logic;
    I2 : in  std_logic;
    I3 : in  std_logic;
    I4 : in  std_logic;
    O  : out std_logic
);
end NX_LUT;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_DFF is
generic (
    dff_edge   : bit       := '0';
    dff_init   : bit       := '0';
    dff_load   : bit       := '0';
    dff_sync   : bit       := '0';
    dff_type   : integer   := 0;
    dff_ctxt   : std_logic := 'U'
);
port (
    I  : in  std_logic;
    CK : in  std_logic;
    L  : in  std_logic;
    R  : in  std_logic;
    O  : out std_logic
);
end NX_DFF;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_BFF is
port (
    I : in  std_logic;
    O : out std_logic
);
end NX_BFF;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_DFR is
generic (
    location   : string  := "";
    iobname    : string  := "";
    path       : integer := 0;
    mode       : integer := 0;
    ring       : integer := 0;
    dff_edge   : bit     := '0';
    dff_init   : bit     := '0';
    dff_load   : bit     := '0';
    dff_sync   : bit     := '0';
    dff_type   : integer := 0
);
port (
    I  : in  std_logic;
    CK : in  std_logic;
    L  : in  std_logic;
    R  : in  std_logic;
    O  : out std_logic
);
end NX_DFR;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_BFR is
generic (
    location   : string := "";
    iobname    : string := "";
    path       : integer := 0;
    mode       : integer := 0;
    data_inv   : bit     := '0';
    ring       : integer := 0
);
port (
    I : in  std_logic;
    O : out std_logic
);
end NX_BFR;

-- =================================================================================================
--   NX_IOB definition                                                                  2017/09/04
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;

entity NX_IOB_I is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  1;
    locked               : bit     := '0'
);
port (
--  I  : in  std_logic;			// To prevent error in instanciation
    C  : in  std_logic;
    T  : in  std_logic;
    IO : in  std_logic;
    O  : out std_logic
);
end NX_IOB_I;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_IOB_O is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  2;
    locked               : bit     := '0'
);
port (
    I  : in  std_logic;
    C  : in  std_logic;
    T  : in  std_logic;
--  O  : out std_logic;			// To prevent error in instanciation
    IO : out std_logic
);
end NX_IOB_O;

----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity NX_IOB is
generic (
    location             : string  := "";
    standard             : string  := "";
    drive                : string  := "";
    differential         : string  := "";
    slewRate             : string  := "";
    termination          : string  := "";
    terminationReference : string  := "";
    turbo                : string  := "";
    weakTermination      : string  := "";
    inputDelayOn         : string  := "";
    inputDelayLine       : string  := "";
    outputDelayOn        : string  := "";
    outputDelayLine      : string  := "";
    inputSignalSlope     : string  := "";
    outputCapacity       : string  := "";
    dynDrive             : string  := "";
    dynInput             : string  := "";
    dynTerm              : string  := "";
    extra                : integer :=  3;
    locked               : bit     := '0'
);
port (
    I  : in    std_logic;
    C  : in    std_logic;
    T  : in    std_logic;
    O  : out   std_logic;
    IO : inout std_logic
);
end NX_IOB;

-- beware following components are only intended for internal use. Do not try to instantiate them.

-- =================================================================================================
--   NX_BUFFER definition                                                               2017/09/11
-- =================================================================================================

-- NX_BUFFER#{{{#
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity NX_BUFFER is
port (
    I : in  std_logic;
    O : out std_logic
);
end NX_BUFFER;
-- #}}}#

-- =================================================================================================
--   NX_CSC definition                                                                  2017/09/26
-- =================================================================================================

-- NX_CSC#{{{#
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity NX_CSC is
port (
    I  : in  std_logic;
    O  : out std_logic
);
end NX_CSC;
-- #}}}#

-- =================================================================================================
--   NX_SCC definition                                                                  2017/09/26
-- =================================================================================================

-- NX_SCC#{{{#
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity NX_SCC is
port (
    I : in  std_logic;
    O : out std_logic
);
end NX_SCC;
-- #}}}#

-- =================================================================================================
--   NX_syn_tp definition                                                               2017/09/11
-- =================================================================================================

-- NX_syn_tp#{{{#
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity NX_syn_tp is
port (
    I : in  std_logic
);
end NX_syn_tp;
-- #}}}#


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity NX_RAM is
generic (
   std_mode     : string := ""; -- standard mode [FAST_2kx18, SLOW_2kx18, NOECNOECC24, ...] empty for raw
   mcka_edge    : bit := '0';   -- 0: rising edge for port A clock - 1: falling edge
   mckb_edge    : bit := '0';   -- 0: rising edge for port B clock - 1: falling edge
   pcka_edge    : bit := '0';   -- 0: rising edge for pipe A clock - 1: falling edge
   pckb_edge    : bit := '0';   -- 0: rising edge for pipe B clock - 1: falling edge
   pipe_ia      : bit := '0';   -- 0: no pipe on port A input  - 1: pipe on port A input
   pipe_ib      : bit := '0';   -- 0: no pipe on port B input  - 1: pipe on port B input
   pipe_oa      : bit := '0';   -- 0: no pipe on port A output - 1: pipe on port A output
   pipe_ob      : bit := '0';   -- 0: no pipe on port B output - 1: pipe on port B output

   raw_config0  : bit_vector( 3 downto 0) := B"0000";			-- PRC
   raw_config1  : bit_vector(15 downto 0) := B"0000000000000000";	-- MOD

   -- For specific NG_LARGE Extended Features
   raw_l_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-LARGE extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_l_extend : bit_vector( 3 downto 0) := B"0000";	    -- Extended modes for NG-LARGE (Scrubbing, test... )

   -- For specific NG_ULTRA Extended Features
   raw_u_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-ULTRA extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_u_extend : bit_vector( 7 downto 0) := B"00000000";   -- Extended modes for NG-ULTRA (Scrubbing, test... )

   mem_ctxt     : string := ""				    -- context initialization
   );
port (
   ACK  : in  std_logic;
   ACKC : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   ACKD : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   ACKR : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   BCK  : in  std_logic;
   BCKC : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   BCKD : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   BCKR : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only

   AI1   : in  std_logic;
   AI2   : in  std_logic;
   AI3   : in  std_logic;
   AI4   : in  std_logic;
   AI5   : in  std_logic;
   AI6   : in  std_logic;
   AI7   : in  std_logic;
   AI8   : in  std_logic;
   AI9   : in  std_logic;
   AI10  : in  std_logic;
   AI11  : in  std_logic;
   AI12  : in  std_logic;
   AI13  : in  std_logic;
   AI14  : in  std_logic;
   AI15  : in  std_logic;
   AI16  : in  std_logic;

   AI17  : in  std_logic;
   AI18  : in  std_logic;
   AI19  : in  std_logic;
   AI20  : in  std_logic;
   AI21  : in  std_logic;
   AI22  : in  std_logic;
   AI23  : in  std_logic;
   AI24  : in  std_logic;

   BI1   : in  std_logic;
   BI2   : in  std_logic;
   BI3   : in  std_logic;
   BI4   : in  std_logic;
   BI5   : in  std_logic;
   BI6   : in  std_logic;
   BI7   : in  std_logic;
   BI8   : in  std_logic;
   BI9   : in  std_logic;
   BI10  : in  std_logic;
   BI11  : in  std_logic;
   BI12  : in  std_logic;
   BI13  : in  std_logic;
   BI14  : in  std_logic;
   BI15  : in  std_logic;
   BI16  : in  std_logic;

   BI17  : in  std_logic;
   BI18  : in  std_logic;
   BI19  : in  std_logic;
   BI20  : in  std_logic;
   BI21  : in  std_logic;
   BI22  : in  std_logic;
   BI23  : in  std_logic;
   BI24  : in  std_logic;

   ACOR  : out std_logic;
   AERR  : out std_logic;
   BCOR  : out std_logic;
   BERR  : out std_logic;

   AO1   : out std_logic;
   AO2   : out std_logic;
   AO3   : out std_logic;
   AO4   : out std_logic;
   AO5   : out std_logic;
   AO6   : out std_logic;
   AO7   : out std_logic;
   AO8   : out std_logic;
   AO9   : out std_logic;
   AO10  : out std_logic;
   AO11  : out std_logic;
   AO12  : out std_logic;
   AO13  : out std_logic;
   AO14  : out std_logic;
   AO15  : out std_logic;
   AO16  : out std_logic;

   AO17  : out std_logic;
   AO18  : out std_logic;
   AO19  : out std_logic;
   AO20  : out std_logic;
   AO21  : out std_logic;
   AO22  : out std_logic;
   AO23  : out std_logic;
   AO24  : out std_logic;

   BO1   : out std_logic;
   BO2   : out std_logic;
   BO3   : out std_logic;
   BO4   : out std_logic;
   BO5   : out std_logic;
   BO6   : out std_logic;
   BO7   : out std_logic;
   BO8   : out std_logic;
   BO9   : out std_logic;
   BO10  : out std_logic;
   BO11  : out std_logic;
   BO12  : out std_logic;
   BO13  : out std_logic;
   BO14  : out std_logic;
   BO15  : out std_logic;
   BO16  : out std_logic;

   BO17  : out std_logic;
   BO18  : out std_logic;
   BO19  : out std_logic;
   BO20  : out std_logic;
   BO21  : out std_logic;
   BO22  : out std_logic;
   BO23  : out std_logic;
   BO24  : out std_logic;

   AA1   : in  std_logic;
   AA2   : in  std_logic;
   AA3   : in  std_logic;
   AA4   : in  std_logic;
   AA5   : in  std_logic;
   AA6   : in  std_logic;

   AA7   : in  std_logic;
   AA8   : in  std_logic;
   AA9   : in  std_logic;
   AA10  : in  std_logic;
   AA11  : in  std_logic;
   AA12  : in  std_logic;
   AA13  : in  std_logic;
   AA14  : in  std_logic;
   AA15  : in  std_logic;
   AA16  : in  std_logic;

   ACS   : in  std_logic;
   AWE   : in  std_logic;
   AR    : in  std_logic;

   BA1   : in  std_logic;
   BA2   : in  std_logic;
   BA3   : in  std_logic;
   BA4   : in  std_logic;
   BA5   : in  std_logic;
   BA6   : in  std_logic;

   BA7   : in  std_logic;
   BA8   : in  std_logic;
   BA9   : in  std_logic;
   BA10  : in  std_logic;
   BA11  : in  std_logic;
   BA12  : in  std_logic;
   BA13  : in  std_logic;
   BA14  : in  std_logic;
   BA15  : in  std_logic;
   BA16  : in  std_logic;

   BCS   : in  std_logic;
   BWE   : in  std_logic;
   BR    : in  std_logic
);
end NX_RAM;

----------------------------------------------------------------------------------------------------

-- =================================================================================================
--   NX_RAM_WRAP definition                                                             2017/09/25
-- =================================================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity NX_RAM_WRAP is
generic (
   std_mode     : string := ""; -- standard mode [FAST_2kx18, SLOW_2kx18, NOECNOECC24, ...] empty for raw
   mcka_edge    : bit := '0';   -- 0: rising edge for port A clock - 1: falling edge
   mckb_edge    : bit := '0';   -- 0: rising edge for port B clock - 1: falling edge
   pcka_edge    : bit := '0';   -- 0: rising edge for pipe A clock - 1: falling edge
   pckb_edge    : bit := '0';   -- 0: rising edge for pipe B clock - 1: falling edge

   pipe_ia      : bit := '0';   -- 0: no pipe on port A input  - 1: pipe on port A input
   pipe_ib      : bit := '0';   -- 0: no pipe on port B input  - 1: pipe on port B input
   pipe_oa      : bit := '0';   -- 0: no pipe on port A output - 1: pipe on port A output
   pipe_ob      : bit := '0';   -- 0: no pipe on port B output - 1: pipe on port B output

   raw_config0  : bit_vector( 3 downto 0) := B"0000";			-- PRC
   raw_config1  : bit_vector(15 downto 0) := B"0000000000000000";	-- MOD

   -- For specific NG_LARGE Extended Features
   raw_l_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-LARGE extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_l_extend : bit_vector( 3 downto 0) := B"0000";	    -- Extended modes for NG-LARGE (Scrubbing, test... )

   -- For specific NG_ULTRA Extended Features
   raw_u_enable : bit := '0';				    -- '0' for NG-MEDIUM, '1' for NG-ULTRA extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_u_extend : bit_vector( 7 downto 0) := B"00000000";   -- Extended modes for NG-ULTRA (Scrubbing, test... )

   mem_ctxt     : string := ""				    -- context initialization
);
port (
   ACK  : in  std_logic;
   ACKD : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   ACKR : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   BCK  : in  std_logic;
   BCKD : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only
   BCKR : in  std_logic;	    -- NG_MEDIUM / NG_LARGE Only

   AI   : in  std_logic_vector(23 downto 0);
   BI   : in  std_logic_vector(23 downto 0);

   ACOR : out std_logic;
   AERR : out std_logic;
   BCOR : out std_logic;
   BERR : out std_logic;

   AO   : out std_logic_vector(23 downto 0);
   BO   : out std_logic_vector(23 downto 0);
   AA   : in  std_logic_vector(15 downto 0);

   ACS  : in  std_logic;
   AWE  : in  std_logic;
   AR   : in  std_logic;

   BA   : in  std_logic_vector(15 downto 0);

   BCS  : in  std_logic;
   BWE  : in  std_logic;
   BR   : in  std_logic
);
end NX_RAM_WRAP;

architecture NX_RTL of NX_RAM_WRAP is
   attribute NX_TYPE :string;
   attribute NX_TYPE of NX_RTL: architecture is "WRAPPER";

component NX_RAM
generic (
   std_mode     : string := ""; -- standard mode [FAST_2kx18, SLOW_2kx18, NOECNOECC24, ...] empty for raw
   mcka_edge    : bit := '0';   -- 0: rising edge for port A clock - 1: falling edge
   mckb_edge    : bit := '0';   -- 0: rising edge for port B clock - 1: falling edge
   pcka_edge    : bit := '0';   -- 0: rising edge for pipe A clock - 1: falling edge
   pckb_edge    : bit := '0';   -- 0: rising edge for pipe B clock - 1: falling edge

   pipe_ia      : bit := '0';   -- 0: no pipe on port A input  - 1: pipe on port A input
   pipe_ib      : bit := '0';   -- 0: no pipe on port B input  - 1: pipe on port B input
   pipe_oa      : bit := '0';   -- 0: no pipe on port A output - 1: pipe on port A output
   pipe_ob      : bit := '0';   -- 0: no pipe on port B output - 1: pipe on port B output

   raw_config0  : bit_vector( 3 downto 0) := B"0000";			-- PRC
   raw_config1  : bit_vector(15 downto 0) := B"0000000000000000";	-- MOD

   raw_l_enable : bit := '0';                         -- '0' for NG-MEDIUM, '1' for NG-LARGE extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_l_extend : bit_vector( 3 downto 0) := B"0000"; -- Extended modes for NG-LARGE (Scrubbing, test... )

   -- For specific NG_ULTRA Extended Features
   raw_u_enable : bit := '0';                         -- '0' for NG-MEDIUM, '1' for NG-ULTRA extended modes (NO_ECC x3 & x6) + scrubbing, test...
   raw_u_extend : bit_vector( 7 downto 0) := B"00000000"; -- Extended modes for NG-ULTRA (Scrubbing, test... )

   mem_ctxt     : string := ""                        -- context initialization
);
port (
   ACK   : in  std_logic;
   ACKC  : in  std_logic;
   ACKD  : in  std_logic;
   ACKR  : in  std_logic;
   BCK   : in  std_logic;
   BCKC  : in  std_logic;
   BCKD  : in  std_logic;
   BCKR  : in  std_logic;

   AI1   : in  std_logic;
   AI2   : in  std_logic;
   AI3   : in  std_logic;
   AI4   : in  std_logic;
   AI5   : in  std_logic;
   AI6   : in  std_logic;
   AI7   : in  std_logic;
   AI8   : in  std_logic;
   AI9   : in  std_logic;
   AI10  : in  std_logic;
   AI11  : in  std_logic;
   AI12  : in  std_logic;
   AI13  : in  std_logic;
   AI14  : in  std_logic;
   AI15  : in  std_logic;
   AI16  : in  std_logic;

   AI17  : in  std_logic;
   AI18  : in  std_logic;
   AI19  : in  std_logic;
   AI20  : in  std_logic;
   AI21  : in  std_logic;
   AI22  : in  std_logic;
   AI23  : in  std_logic;
   AI24  : in  std_logic;

   BI1   : in  std_logic;
   BI2   : in  std_logic;
   BI3   : in  std_logic;
   BI4   : in  std_logic;
   BI5   : in  std_logic;
   BI6   : in  std_logic;
   BI7   : in  std_logic;
   BI8   : in  std_logic;
   BI9   : in  std_logic;
   BI10  : in  std_logic;
   BI11  : in  std_logic;
   BI12  : in  std_logic;
   BI13  : in  std_logic;
   BI14  : in  std_logic;
   BI15  : in  std_logic;
   BI16  : in  std_logic;

   BI17  : in  std_logic;
   BI18  : in  std_logic;
   BI19  : in  std_logic;
   BI20  : in  std_logic;
   BI21  : in  std_logic;
   BI22  : in  std_logic;
   BI23  : in  std_logic;
   BI24  : in  std_logic;

   ACOR  : out std_logic;
   AERR  : out std_logic;
   BCOR  : out std_logic;
   BERR  : out std_logic;

   AO1   : out std_logic;
   AO2   : out std_logic;
   AO3   : out std_logic;
   AO4   : out std_logic;
   AO5   : out std_logic;
   AO6   : out std_logic;
   AO7   : out std_logic;
   AO8   : out std_logic;
   AO9   : out std_logic;
   AO10  : out std_logic;
   AO11  : out std_logic;
   AO12  : out std_logic;
   AO13  : out std_logic;
   AO14  : out std_logic;
   AO15  : out std_logic;
   AO16  : out std_logic;

   AO17  : out std_logic;
   AO18  : out std_logic;
   AO19  : out std_logic;
   AO20  : out std_logic;
   AO21  : out std_logic;
   AO22  : out std_logic;
   AO23  : out std_logic;
   AO24  : out std_logic;

   BO1   : out std_logic;
   BO2   : out std_logic;
   BO3   : out std_logic;
   BO4   : out std_logic;
   BO5   : out std_logic;
   BO6   : out std_logic;
   BO7   : out std_logic;
   BO8   : out std_logic;
   BO9   : out std_logic;
   BO10  : out std_logic;
   BO11  : out std_logic;
   BO12  : out std_logic;
   BO13  : out std_logic;
   BO14  : out std_logic;
   BO15  : out std_logic;
   BO16  : out std_logic;

   BO17  : out std_logic;
   BO18  : out std_logic;
   BO19  : out std_logic;
   BO20  : out std_logic;
   BO21  : out std_logic;
   BO22  : out std_logic;
   BO23  : out std_logic;
   BO24  : out std_logic;

   AA1   : in  std_logic;
   AA2   : in  std_logic;
   AA3   : in  std_logic;
   AA4   : in  std_logic;
   AA5   : in  std_logic;
   AA6   : in  std_logic;

   AA7   : in  std_logic;
   AA8   : in  std_logic;
   AA9   : in  std_logic;
   AA10  : in  std_logic;
   AA11  : in  std_logic;
   AA12  : in  std_logic;
   AA13  : in  std_logic;
   AA14  : in  std_logic;
   AA15  : in  std_logic;
   AA16  : in  std_logic;

   ACS   : in  std_logic;
   AWE   : in  std_logic;
   AR    : in  std_logic;

   BA1   : in  std_logic;
   BA2   : in  std_logic;
   BA3   : in  std_logic;
   BA4   : in  std_logic;
   BA5   : in  std_logic;
   BA6   : in  std_logic;

   BA7   : in  std_logic;
   BA8   : in  std_logic;
   BA9   : in  std_logic;
   BA10  : in  std_logic;
   BA11  : in  std_logic;
   BA12  : in  std_logic;
   BA13  : in  std_logic;
   BA14  : in  std_logic;
   BA15  : in  std_logic;
   BA16  : in  std_logic;

   BCS   : in  std_logic;
   BWE   : in  std_logic;
   BR    : in  std_logic
);
end component;

begin

ram: NX_RAM generic map (
   std_mode     => std_mode,
   mcka_edge    => mcka_edge,
   mckb_edge    => mckb_edge,
   pcka_edge    => pcka_edge,
   pckb_edge    => pckb_edge,
   pipe_ia      => pipe_ia,
   pipe_ib      => pipe_ib,
   pipe_oa      => pipe_oa,
   pipe_ob      => pipe_ob,
   raw_config0  => raw_config0,
   raw_config1  => raw_config1,
   raw_l_enable => raw_l_enable,
   raw_u_enable => raw_u_enable,
   raw_l_extend => raw_l_extend,
   raw_u_extend => raw_u_extend,
   mem_ctxt     => mem_ctxt
)
port map(
   ACK   => ACK,
   ACKC  => ACK,
   ACKD  => ACKD,
   ACKR  => ACKR,
   BCK   => BCK,
   BCKC  => BCK,
   BCKD  => BCKD,
   BCKR  => BCKR,

   AI1   => AI(0),
   AI2   => AI(1),
   AI3   => AI(2),
   AI4   => AI(3),
   AI5   => AI(4),
   AI6   => AI(5),
   AI7   => AI(6),
   AI8   => AI(7),
   AI9   => AI(8),
   AI10  => AI(9),
   AI11  => AI(10),
   AI12  => AI(11),
   AI13  => AI(12),
   AI14  => AI(13),
   AI15  => AI(14),
   AI16  => AI(15),

   AI17  => AI(16),
   AI18  => AI(17),
   AI19  => AI(18),
   AI20  => AI(19),
   AI21  => AI(20),
   AI22  => AI(21),
   AI23  => AI(22),
   AI24  => AI(23),

   BI1   => BI(0),
   BI2   => BI(1),
   BI3   => BI(2),
   BI4   => BI(3),
   BI5   => BI(4),
   BI6   => BI(5),
   BI7   => BI(6),
   BI8   => BI(7),
   BI9   => BI(8),
   BI10  => BI(9),
   BI11  => BI(10),
   BI12  => BI(11),
   BI13  => BI(12),
   BI14  => BI(13),
   BI15  => BI(14),
   BI16  => BI(15),

   BI17  => BI(16),
   BI18  => BI(17),
   BI19  => BI(18),
   BI20  => BI(19),
   BI21  => BI(20),
   BI22  => BI(21),
   BI23  => BI(22),
   BI24  => BI(23),

   ACOR  => ACOR,
   AERR  => AERR,
   BCOR  => BCOR,
   BERR  => BERR,

   AO1   => AO(0),
   AO2   => AO(1),
   AO3   => AO(2),
   AO4   => AO(3),
   AO5   => AO(4),
   AO6   => AO(5),
   AO7   => AO(6),
   AO8   => AO(7),
   AO9   => AO(8),
   AO10  => AO(9),
   AO11  => AO(10),
   AO12  => AO(11),
   AO13  => AO(12),
   AO14  => AO(13),
   AO15  => AO(14),
   AO16  => AO(15),

   AO17  => AO(16),
   AO18  => AO(17),
   AO19  => AO(18),
   AO20  => AO(19),
   AO21  => AO(20),
   AO22  => AO(21),
   AO23  => AO(22),
   AO24  => AO(23),

   BO1   => BO(0),
   BO2   => BO(1),
   BO3   => BO(2),
   BO4   => BO(3),
   BO5   => BO(4),
   BO6   => BO(5),
   BO7   => BO(6),
   BO8   => BO(7),
   BO9   => BO(8),
   BO10  => BO(9),
   BO11  => BO(10),
   BO12  => BO(11),
   BO13  => BO(12),
   BO14  => BO(13),
   BO15  => BO(14),
   BO16  => BO(15),

   BO17  => BO(16),
   BO18  => BO(17),
   BO19  => BO(18),
   BO20  => BO(19),
   BO21  => BO(20),
   BO22  => BO(21),
   BO23  => BO(22),
   BO24  => BO(23),

   AA1   => AA(0),
   AA2   => AA(1),
   AA3   => AA(2),
   AA4   => AA(3),
   AA5   => AA(4),
   AA6   => AA(5),

   AA7   => AA(6),
   AA8   => AA(7),
   AA9   => AA(8),
   AA10  => AA(9),
   AA11  => AA(10),
   AA12  => AA(11),
   AA13  => AA(12),
   AA14  => AA(13),
   AA15  => AA(14),
   AA16  => AA(15),

   ACS   => ACS,
   AWE   => AWE,
   AR    => AR,

   BA1   => BA(0),
   BA2   => BA(1),
   BA3   => BA(2),
   BA4   => BA(3),
   BA5   => BA(4),
   BA6   => BA(5),

   BA7   => BA(6),
   BA8   => BA(7),
   BA9   => BA(8),
   BA10  => BA(9),
   BA11  => BA(10),
   BA12  => BA(11),
   BA13  => BA(12),
   BA14  => BA(13),
   BA15  => BA(14),
   BA16  => BA(15),

   BCS   => BCS,
   BWE   => BWE,
   BR    => BR
   );

end NX_RTL;
architecture NX_RTL of NX_CDC_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CDC_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_CDC_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_FIFO_CDC_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CDC_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (XRCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_CDC_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_DSP_L_BOX is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "BOX";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DSP_L_BOX";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_DSP_L_BOX doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_RAM_L_BOX is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "BOX";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RAM_L_BOX";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (ACK) begin				    -- Dummy input for syntax analysis
	report "Model NX_RAM_L_BOX doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_DSP_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DSP_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_DSP_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_DSP is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DSP";
begin

fail : if NX_SYMBOL /= "NG_M" generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_DSP doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_DSP_U_BOX is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "BOX";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DSP_U_BOX";
begin

fail : if (NX_SYMBOL /= "NG_U") and (NX_SYMBOL /= "NG_C") generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_DSP_U_BOX doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;


end NX_RTL;
architecture NX_RTL of NX_RAM_U_BOX is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "BOX";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RAM_U_BOX";
begin

fail : if (NX_SYMBOL /= "NG_U") and (NX_SYMBOL /= "NG_C") generate
    process (ACK) begin				    -- Dummy input for syntax analysis
	report "Model NX_RAM_U_BOX doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_DSP_U is
    attribute NX_TYPE           : string;
    attribute NX_TYPE of NX_RTL : architecture is "PHY";

    attribute NX_USE            : string;
    attribute NX_USE of NX_RTL  : architecture is "NX_DSP_U";
begin

fail : if (NX_SYMBOL /= "NG_U") and (NX_SYMBOL /= "NG_C") generate
    process (CK) begin				    -- Dummy input for syntax analysis
	report "Model NX_DSP_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_FIFO_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_FIFO_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (RCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_FIFO_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_GCK_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_GCK_U";

begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (SI1) begin				    -- Dummy input for syntax analysis
	report "Model NX_GCK_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_CRX_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CRX_L";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (RX_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_CRX_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_CTX_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CTX_L";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CLK_E_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_CTX_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_PMA_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_PMA_L";
    attribute NX_USE of LINK_TX0: signal is "LINK";
    attribute NX_USE of LINK_TX1: signal is "LINK";
    attribute NX_USE of LINK_TX2: signal is "LINK";
    attribute NX_USE of LINK_TX3: signal is "LINK";
    attribute NX_USE of LINK_TX4: signal is "LINK";
    attribute NX_USE of LINK_TX5: signal is "LINK";
    attribute NX_USE of LINK_RX0: signal is "LINK";
    attribute NX_USE of LINK_RX1: signal is "LINK";
    attribute NX_USE of LINK_RX2: signal is "LINK";
    attribute NX_USE of LINK_RX3: signal is "LINK";
    attribute NX_USE of LINK_RX4: signal is "LINK";
    attribute NX_USE of LINK_RX5: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CLK_REF_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_PMA_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_CRX_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CRX_U";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (RST_N_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_CRX_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_CTX_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CTX_U";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CLK_E_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_CTX_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_PMA_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_PMA_U";
    attribute NX_USE of LINK_TX0: signal is "LINK";
    attribute NX_USE of LINK_TX1: signal is "LINK";
    attribute NX_USE of LINK_TX2: signal is "LINK";
    attribute NX_USE of LINK_TX3: signal is "LINK";
    attribute NX_USE of LINK_RX0: signal is "LINK";
    attribute NX_USE of LINK_RX1: signal is "LINK";
    attribute NX_USE of LINK_RX2: signal is "LINK";
    attribute NX_USE of LINK_RX3: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CLK_REF_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_PMA_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_IOM_L is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;


architecture NX_RTL of NX_IOM_CONTROL_L is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_CONTROL_L";
    attribute NX_USE of LINK1  : signal is "LINK";
    attribute NX_USE of LINK2  : signal is "LINK";
    attribute NX_USE of LINK3  : signal is "LINK";
    attribute NX_USE of LINK4  : signal is "LINK";
    attribute NX_USE of LINK5  : signal is "LINK";
    attribute NX_USE of LINK6  : signal is "LINK";
    attribute NX_USE of LINK7  : signal is "LINK";
    attribute NX_USE of LINK8  : signal is "LINK";
    attribute NX_USE of LINK9  : signal is "LINK";
    attribute NX_USE of LINK10 : signal is "LINK";
    attribute NX_USE of LINK11 : signal is "LINK";
    attribute NX_USE of LINK12 : signal is "LINK";
    attribute NX_USE of LINK13 : signal is "LINK";
    attribute NX_USE of LINK14 : signal is "LINK";
    attribute NX_USE of LINK15 : signal is "LINK";
    attribute NX_USE of LINK16 : signal is "LINK";
    attribute NX_USE of LINK17 : signal is "LINK";
    attribute NX_USE of LINK18 : signal is "LINK";
    attribute NX_USE of LINK19 : signal is "LINK";
    attribute NX_USE of LINK20 : signal is "LINK";
    attribute NX_USE of LINK21 : signal is "LINK";
    attribute NX_USE of LINK22 : signal is "LINK";
    attribute NX_USE of LINK23 : signal is "LINK";
    attribute NX_USE of LINK24 : signal is "LINK";
    attribute NX_USE of LINK25 : signal is "LINK";
    attribute NX_USE of LINK26 : signal is "LINK";
    attribute NX_USE of LINK27 : signal is "LINK";
    attribute NX_USE of LINK28 : signal is "LINK";
    attribute NX_USE of LINK29 : signal is "LINK";
    attribute NX_USE of LINK30 : signal is "LINK";
    attribute NX_USE of LINK31 : signal is "LINK";
    attribute NX_USE of LINK32 : signal is "LINK";
    attribute NX_USE of LINK33 : signal is "LINK";
    attribute NX_USE of LINK34 : signal is "LINK";

begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_CONTROL_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_IOM_DRIVER_M is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_DRIVER_M";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_M" and NX_SYMBOL /= "NG_L" generate
    process (CTI) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_DRIVER_M doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_IOM_SERDES_M is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_SERDES_M";
    attribute NX_USE of LINKP: signal is "LINK";
    attribute NX_USE of LINKN: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_M" and NX_SYMBOL /= "NG_L" generate
    process (RTCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_SERDES_M doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_IOM is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM";
begin

fail : if NX_SYMBOL /= "NG_M" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_IOM_CONTROL_M is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_CONTROL_M";
    attribute NX_USE of LINK1  : signal is "LINK";
    attribute NX_USE of LINK2  : signal is "LINK";
    attribute NX_USE of LINK3  : signal is "LINK";
    attribute NX_USE of LINK4  : signal is "LINK";
    attribute NX_USE of LINK5  : signal is "LINK";
    attribute NX_USE of LINK6  : signal is "LINK";
    attribute NX_USE of LINK7  : signal is "LINK";
    attribute NX_USE of LINK8  : signal is "LINK";
    attribute NX_USE of LINK9  : signal is "LINK";
    attribute NX_USE of LINK10 : signal is "LINK";
    attribute NX_USE of LINK11 : signal is "LINK";
    attribute NX_USE of LINK12 : signal is "LINK";
    attribute NX_USE of LINK13 : signal is "LINK";
    attribute NX_USE of LINK14 : signal is "LINK";
    attribute NX_USE of LINK15 : signal is "LINK";
    attribute NX_USE of LINK16 : signal is "LINK";
    attribute NX_USE of LINK17 : signal is "LINK";
    attribute NX_USE of LINK18 : signal is "LINK";
    attribute NX_USE of LINK19 : signal is "LINK";
    attribute NX_USE of LINK20 : signal is "LINK";
    attribute NX_USE of LINK21 : signal is "LINK";
    attribute NX_USE of LINK22 : signal is "LINK";
    attribute NX_USE of LINK23 : signal is "LINK";
    attribute NX_USE of LINK24 : signal is "LINK";
    attribute NX_USE of LINK25 : signal is "LINK";
    attribute NX_USE of LINK26 : signal is "LINK";
    attribute NX_USE of LINK27 : signal is "LINK";
    attribute NX_USE of LINK28 : signal is "LINK";
    attribute NX_USE of LINK29 : signal is "LINK";
    attribute NX_USE of LINK30 : signal is "LINK";
    attribute NX_USE of LINK31 : signal is "LINK";
    attribute NX_USE of LINK32 : signal is "LINK";
    attribute NX_USE of LINK33 : signal is "LINK";
    attribute NX_USE of LINK34 : signal is "LINK";

begin

fail : if NX_SYMBOL /= "NG_M" and NX_SYMBOL /= "NG_L" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_CONTROL_M doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;
end NX_RTL;
architecture NX_RTL of NX_IOM_DRIVER_U is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_DRIVER_U";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CTI) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_DRIVER_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_IOM_SERDES_U is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_SERDES_U";
    attribute NX_USE of LINK: signal is "LINK";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (FCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_SERDES_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_IOM_U is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;


architecture NX_RTL of NX_IOM_CONTROL_U is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOM_CONTROL_U";
    attribute NX_USE of LINK1  : signal is "LINK";
    attribute NX_USE of LINK2  : signal is "LINK";
    attribute NX_USE of LINK3  : signal is "LINK";
    attribute NX_USE of LINK4  : signal is "LINK";
    attribute NX_USE of LINK5  : signal is "LINK";
    attribute NX_USE of LINK6  : signal is "LINK";
    attribute NX_USE of LINK7  : signal is "LINK";
    attribute NX_USE of LINK8  : signal is "LINK";
    attribute NX_USE of LINK9  : signal is "LINK";
    attribute NX_USE of LINK10 : signal is "LINK";
    attribute NX_USE of LINK11 : signal is "LINK";
    attribute NX_USE of LINK12 : signal is "LINK";
    attribute NX_USE of LINK13 : signal is "LINK";
    attribute NX_USE of LINK14 : signal is "LINK";
    attribute NX_USE of LINK15 : signal is "LINK";
    attribute NX_USE of LINK16 : signal is "LINK";
    attribute NX_USE of LINK17 : signal is "LINK";
    attribute NX_USE of LINK18 : signal is "LINK";
    attribute NX_USE of LINK19 : signal is "LINK";
    attribute NX_USE of LINK20 : signal is "LINK";
    attribute NX_USE of LINK21 : signal is "LINK";
    attribute NX_USE of LINK22 : signal is "LINK";
    attribute NX_USE of LINK23 : signal is "LINK";
    attribute NX_USE of LINK24 : signal is "LINK";
    attribute NX_USE of LINK25 : signal is "LINK";
    attribute NX_USE of LINK26 : signal is "LINK";
    attribute NX_USE of LINK27 : signal is "LINK";
    attribute NX_USE of LINK28 : signal is "LINK";
    attribute NX_USE of LINK29 : signal is "LINK";
    attribute NX_USE of LINK30 : signal is "LINK";
    attribute NX_USE of LINK31 : signal is "LINK";
    attribute NX_USE of LINK32 : signal is "LINK";
    attribute NX_USE of LINK33 : signal is "LINK";
    attribute NX_USE of LINK34 : signal is "LINK";

begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_IOM_CONTROL_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
-- =================================================================================================
--   NX_PLL_L definition                                                                2018/11/30
-- =================================================================================================

architecture NX_RTL of NX_PLL_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_PLL_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (REF) begin				    -- Dummy input for syntax analysis
	report "Model NX_PLL_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

-- =================================================================================================
--   NX_WFG_L definition                                                                2018/11/30
-- =================================================================================================

architecture NX_RTL of NX_WFG_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_WFG_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (SI) begin				    -- Dummy input for syntax analysis
	report "Model NX_WFG_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

-- =================================================================================================
--   NX_PLL definition                                                                  2017/09/19
-- =================================================================================================

architecture NX_RTL of NX_PLL is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_PLL";
begin

fail : if NX_SYMBOL /= "NG_M" generate
    process (REF) begin				    -- Dummy input for syntax analysis
	report "Model NX_PLL doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

-- =================================================================================================
--   NX_WFG definition                                                                  2017/09/19
-- =================================================================================================

architecture NX_RTL of NX_WFG is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_WFG";
begin

fail : if NX_SYMBOL /= "NG_M" generate
    process (SI) begin				    -- Dummy input for syntax analysis
	report "Model NX_WFG doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_PLL_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_PLL_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (REF) begin				    -- Dummy input for syntax analysis
	report "Model NX_PLL_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_WFG_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_WFG_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (R) begin				    -- Dummy input for syntax analysis
	report "Model NX_WFG_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_R5_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_R5_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (CK_I) begin				    -- Dummy input for syntax analysis
	report "Model NX_R5_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_RB is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RB";
begin

fail : if NX_SYMBOL /= "NG_C" generate
    process (CK1) begin				    -- Dummy input for syntax analysis
	report "Model NX_RB doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_RFB_L is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RFB_L";
begin

fail : if NX_SYMBOL /= "NG_L" generate
    process (RCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_RFB_L doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
-- =================================================================================================
--   NX_RFB_M definition                                                                 2017/09/19
-- =================================================================================================

architecture NX_RTL of NX_RFB_M is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RFB_M";
begin

fail : if NX_SYMBOL /= "NG_M" generate
    process (WCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_RFB_M doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;

architecture NX_RTL of NX_CKS is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CKS";
begin

fail : if (NX_SYMBOL /= "NG_M") and (NX_SYMBOL /= "NG_L") generate
    process (CKI) begin				    -- Dummy input for syntax analysis
	report "Model NX_CKS doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_CDC_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CDC_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (CK1) begin				    -- Dummy input for syntax analysis
	report "Model NX_CDC_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_RFB_U is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RFB_U";
begin

fail : if NX_SYMBOL /= "NG_U" and NX_SYMBOL /= "NG_C" generate
    process (WCK) begin				    -- Dummy input for syntax analysis
	report "Model NX_RFB_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_SERVICE_U is
attribute NX_TYPE :string;
attribute NX_TYPE of NX_RTL: architecture is "PHY";

attribute NX_USE :string;
attribute NX_USE of NX_RTL: architecture is "NX_SERVICE_U";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (fabric_otp_user_tst_scanenable_i) begin				    -- Dummy input for syntax analysis
	report "Model NX_SERVICE_U doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
architecture NX_RTL of NX_SOC_INTERFACE is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_SOC_INTERFACE";
begin

fail : if NX_SYMBOL /= "NG_U" generate
    process (fabric_lowskew_o1) begin				    -- Dummy input for syntax analysis
	report "Model NX_SOC_INTERFACE doesn't belong to " & NX_FAMILY & " family" severity error;
    end process;
end generate;

end NX_RTL;
-- =================================================================================================
--   NX_BD definition                                                                   2018/06/19
-- =================================================================================================

architecture NX_RTL of NX_BD is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_BD";
begin
end NX_RTL;

-- =================================================================================================
--   NX_CY definition                                                                   2017/09/19
-- =================================================================================================

architecture NX_RTL of NX_CY is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_CY";
begin
end NX_RTL;

architecture NX_RTL of NX_ECC is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_ECC";
begin
end NX_RTL;
-- =================================================================================================
--   NX_LUT definition                                                                  2017/09/04
-- =================================================================================================

architecture NX_RTL of NX_LUT is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_LUT";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_DFF is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DFF";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_BFF is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_BFF";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_DFR is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_DFR";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_BFR is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_BFR";
begin
end NX_RTL;

-- =================================================================================================
--   NX_IOB definition                                                                  2017/09/04
-- =================================================================================================

architecture NX_RTL of NX_IOB_I is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOB";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_IOB_O is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOB";
begin
end NX_RTL;

----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_IOB is
    attribute NX_TYPE: string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE: string;
    attribute NX_USE of NX_RTL: architecture is "NX_IOB";
begin
end NX_RTL;

-- =================================================================================================
--   NX_syn_tp definition                                                               2017/09/11
-- =================================================================================================

-- NX_syn_tp#
----------------------------------------------------------------------------------------------------

architecture NX_RTL of NX_syn_tp is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_syn_tp";
begin
end NX_RTL;

-- =================================================================================================
--   NX_RAM definition                                                                  2017/09/25
-- =================================================================================================

architecture NX_RTL of NX_RAM is
    attribute NX_TYPE :string;
    attribute NX_TYPE of NX_RTL: architecture is "PHY";

    attribute NX_USE :string;
    attribute NX_USE of NX_RTL: architecture is "NX_RAM";
begin
end NX_RTL;
