--
-- VHDL Architecture Bachelor.counter_to_aqu.test
--
-- Created:
--          by - christop.grobety.UNKNOWN (WE2332207)
--          at - 13:54:32 30.05.2023
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE test OF counter_to_aqu IS
BEGIN
END ARCHITECTURE test;

