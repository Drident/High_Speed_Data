architecture studentVersion of interpolatorTrigger is

begin

  triggerOut <= '0';

end studentVersion;
