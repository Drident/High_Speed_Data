--
-- VHDL Architecture Bachelor.ADC_Write.STUDENT_VTEST
--
-- Created:
--          by - christop.grobety.UNKNOWN (WE2332207)
--          at - 11:47:26 28.06.2023
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE STUDENT_VTEST OF ADC_Write IS
BEGIN
END ARCHITECTURE STUDENT_VTEST;

