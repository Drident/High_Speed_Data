--
-- VHDL Architecture Bachelor.mux_test.test
--
-- Created:
--          by - christop.grobety.UNKNOWN (WE2332207)
--          at - 13:15:49 30.05.2023
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE test OF mux_test IS
BEGIN
END ARCHITECTURE test;

